/*******************************************************************************
  Copyright 2019 Xi'an Jiaotong University

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
*******************************************************************************/

module xpb_16_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000100000000000000000000000000000000ffffffff0000000000000001;
		5'b00010:	xpb = 256'h0000000200000000000000000000000000000001fffffffe0000000000000002;
		5'b00011:	xpb = 256'h0000000300000000000000000000000000000002fffffffd0000000000000003;
		5'b00100:	xpb = 256'h0000000400000000000000000000000000000003fffffffc0000000000000004;
		5'b00101:	xpb = 256'h0000000500000000000000000000000000000004fffffffb0000000000000005;
		5'b00110:	xpb = 256'h0000000600000000000000000000000000000005fffffffa0000000000000006;
		5'b00111:	xpb = 256'h0000000700000000000000000000000000000006fffffff90000000000000007;
		5'b01000:	xpb = 256'h0000000800000000000000000000000000000007fffffff80000000000000008;
		5'b01001:	xpb = 256'h0000000900000000000000000000000000000008fffffff70000000000000009;
		5'b01010:	xpb = 256'h0000000a00000000000000000000000000000009fffffff6000000000000000a;
		5'b01011:	xpb = 256'h0000000b0000000000000000000000000000000afffffff5000000000000000b;
		5'b01100:	xpb = 256'h0000000c0000000000000000000000000000000bfffffff4000000000000000c;
		5'b01101:	xpb = 256'h0000000d0000000000000000000000000000000cfffffff3000000000000000d;
		5'b01110:	xpb = 256'h0000000e0000000000000000000000000000000dfffffff2000000000000000e;
		5'b01111:	xpb = 256'h0000000f0000000000000000000000000000000efffffff1000000000000000f;
		5'b10000:	xpb = 256'h000000100000000000000000000000000000000ffffffff00000000000000010;
		5'b10001:	xpb = 256'h0000001100000000000000000000000000000010ffffffef0000000000000011;
		5'b10010:	xpb = 256'h0000001200000000000000000000000000000011ffffffee0000000000000012;
		5'b10011:	xpb = 256'h0000001300000000000000000000000000000012ffffffed0000000000000013;
		5'b10100:	xpb = 256'h0000001400000000000000000000000000000013ffffffec0000000000000014;
		5'b10101:	xpb = 256'h0000001500000000000000000000000000000014ffffffeb0000000000000015;
		5'b10110:	xpb = 256'h0000001600000000000000000000000000000015ffffffea0000000000000016;
		5'b10111:	xpb = 256'h0000001700000000000000000000000000000016ffffffe90000000000000017;
		5'b11000:	xpb = 256'h0000001800000000000000000000000000000017ffffffe80000000000000018;
		5'b11001:	xpb = 256'h0000001900000000000000000000000000000018ffffffe70000000000000019;
		5'b11010:	xpb = 256'h0000001a00000000000000000000000000000019ffffffe6000000000000001a;
		5'b11011:	xpb = 256'h0000001b0000000000000000000000000000001affffffe5000000000000001b;
		5'b11100:	xpb = 256'h0000001c0000000000000000000000000000001bffffffe4000000000000001c;
		5'b11101:	xpb = 256'h0000001d0000000000000000000000000000001cffffffe3000000000000001d;
		5'b11110:	xpb = 256'h0000001e0000000000000000000000000000001dffffffe2000000000000001e;
		5'b11111:	xpb = 256'h0000001f0000000000000000000000000000001effffffe1000000000000001f;
	endcase
end
endmodule

module xpb_16_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h000000200000000000000000000000000000001fffffffe00000000000000020;
		6'b000010:	xpb = 256'h000000400000000000000000000000000000003fffffffc00000000000000040;
		6'b000011:	xpb = 256'h000000600000000000000000000000000000005fffffffa00000000000000060;
		6'b000100:	xpb = 256'h000000800000000000000000000000000000007fffffff800000000000000080;
		6'b000101:	xpb = 256'h000000a00000000000000000000000000000009fffffff6000000000000000a0;
		6'b000110:	xpb = 256'h000000c0000000000000000000000000000000bfffffff4000000000000000c0;
		6'b000111:	xpb = 256'h000000e0000000000000000000000000000000dfffffff2000000000000000e0;
		6'b001000:	xpb = 256'h00000100000000000000000000000000000000ffffffff000000000000000100;
		6'b001001:	xpb = 256'h000001200000000000000000000000000000011ffffffee00000000000000120;
		6'b001010:	xpb = 256'h000001400000000000000000000000000000013ffffffec00000000000000140;
		6'b001011:	xpb = 256'h000001600000000000000000000000000000015ffffffea00000000000000160;
		6'b001100:	xpb = 256'h000001800000000000000000000000000000017ffffffe800000000000000180;
		6'b001101:	xpb = 256'h000001a00000000000000000000000000000019ffffffe6000000000000001a0;
		6'b001110:	xpb = 256'h000001c0000000000000000000000000000001bffffffe4000000000000001c0;
		6'b001111:	xpb = 256'h000001e0000000000000000000000000000001dffffffe2000000000000001e0;
		6'b010000:	xpb = 256'h00000200000000000000000000000000000001fffffffe000000000000000200;
		6'b010001:	xpb = 256'h000002200000000000000000000000000000021ffffffde00000000000000220;
		6'b010010:	xpb = 256'h000002400000000000000000000000000000023ffffffdc00000000000000240;
		6'b010011:	xpb = 256'h000002600000000000000000000000000000025ffffffda00000000000000260;
		6'b010100:	xpb = 256'h000002800000000000000000000000000000027ffffffd800000000000000280;
		6'b010101:	xpb = 256'h000002a00000000000000000000000000000029ffffffd6000000000000002a0;
		6'b010110:	xpb = 256'h000002c0000000000000000000000000000002bffffffd4000000000000002c0;
		6'b010111:	xpb = 256'h000002e0000000000000000000000000000002dffffffd2000000000000002e0;
		6'b011000:	xpb = 256'h00000300000000000000000000000000000002fffffffd000000000000000300;
		6'b011001:	xpb = 256'h000003200000000000000000000000000000031ffffffce00000000000000320;
		6'b011010:	xpb = 256'h000003400000000000000000000000000000033ffffffcc00000000000000340;
		6'b011011:	xpb = 256'h000003600000000000000000000000000000035ffffffca00000000000000360;
		6'b011100:	xpb = 256'h000003800000000000000000000000000000037ffffffc800000000000000380;
		6'b011101:	xpb = 256'h000003a00000000000000000000000000000039ffffffc6000000000000003a0;
		6'b011110:	xpb = 256'h000003c0000000000000000000000000000003bffffffc4000000000000003c0;
		6'b011111:	xpb = 256'h000003e0000000000000000000000000000003dffffffc2000000000000003e0;
		6'b100000:	xpb = 256'h00000400000000000000000000000000000003fffffffc000000000000000400;
		6'b100001:	xpb = 256'h000004200000000000000000000000000000041ffffffbe00000000000000420;
		6'b100010:	xpb = 256'h000004400000000000000000000000000000043ffffffbc00000000000000440;
		6'b100011:	xpb = 256'h000004600000000000000000000000000000045ffffffba00000000000000460;
		6'b100100:	xpb = 256'h000004800000000000000000000000000000047ffffffb800000000000000480;
		6'b100101:	xpb = 256'h000004a00000000000000000000000000000049ffffffb6000000000000004a0;
		6'b100110:	xpb = 256'h000004c0000000000000000000000000000004bffffffb4000000000000004c0;
		6'b100111:	xpb = 256'h000004e0000000000000000000000000000004dffffffb2000000000000004e0;
		6'b101000:	xpb = 256'h00000500000000000000000000000000000004fffffffb000000000000000500;
		6'b101001:	xpb = 256'h000005200000000000000000000000000000051ffffffae00000000000000520;
		6'b101010:	xpb = 256'h000005400000000000000000000000000000053ffffffac00000000000000540;
		6'b101011:	xpb = 256'h000005600000000000000000000000000000055ffffffaa00000000000000560;
		6'b101100:	xpb = 256'h000005800000000000000000000000000000057ffffffa800000000000000580;
		6'b101101:	xpb = 256'h000005a00000000000000000000000000000059ffffffa6000000000000005a0;
		6'b101110:	xpb = 256'h000005c0000000000000000000000000000005bffffffa4000000000000005c0;
		6'b101111:	xpb = 256'h000005e0000000000000000000000000000005dffffffa2000000000000005e0;
		6'b110000:	xpb = 256'h00000600000000000000000000000000000005fffffffa000000000000000600;
		6'b110001:	xpb = 256'h000006200000000000000000000000000000061ffffff9e00000000000000620;
		6'b110010:	xpb = 256'h000006400000000000000000000000000000063ffffff9c00000000000000640;
		6'b110011:	xpb = 256'h000006600000000000000000000000000000065ffffff9a00000000000000660;
		6'b110100:	xpb = 256'h000006800000000000000000000000000000067ffffff9800000000000000680;
		6'b110101:	xpb = 256'h000006a00000000000000000000000000000069ffffff96000000000000006a0;
		6'b110110:	xpb = 256'h000006c0000000000000000000000000000006bffffff94000000000000006c0;
		6'b110111:	xpb = 256'h000006e0000000000000000000000000000006dffffff92000000000000006e0;
		6'b111000:	xpb = 256'h00000700000000000000000000000000000006fffffff9000000000000000700;
		6'b111001:	xpb = 256'h000007200000000000000000000000000000071ffffff8e00000000000000720;
		6'b111010:	xpb = 256'h000007400000000000000000000000000000073ffffff8c00000000000000740;
		6'b111011:	xpb = 256'h000007600000000000000000000000000000075ffffff8a00000000000000760;
		6'b111100:	xpb = 256'h000007800000000000000000000000000000077ffffff8800000000000000780;
		6'b111101:	xpb = 256'h000007a00000000000000000000000000000079ffffff86000000000000007a0;
		6'b111110:	xpb = 256'h000007c0000000000000000000000000000007bffffff84000000000000007c0;
		6'b111111:	xpb = 256'h000007e0000000000000000000000000000007dffffff82000000000000007e0;
	endcase
end
endmodule

module xpb_16_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00000800000000000000000000000000000007fffffff8000000000000000800;
		6'b000010:	xpb = 256'h0000100000000000000000000000000000000ffffffff0000000000000001000;
		6'b000011:	xpb = 256'h00001800000000000000000000000000000017ffffffe8000000000000001800;
		6'b000100:	xpb = 256'h0000200000000000000000000000000000001fffffffe0000000000000002000;
		6'b000101:	xpb = 256'h00002800000000000000000000000000000027ffffffd8000000000000002800;
		6'b000110:	xpb = 256'h0000300000000000000000000000000000002fffffffd0000000000000003000;
		6'b000111:	xpb = 256'h00003800000000000000000000000000000037ffffffc8000000000000003800;
		6'b001000:	xpb = 256'h0000400000000000000000000000000000003fffffffc0000000000000004000;
		6'b001001:	xpb = 256'h00004800000000000000000000000000000047ffffffb8000000000000004800;
		6'b001010:	xpb = 256'h0000500000000000000000000000000000004fffffffb0000000000000005000;
		6'b001011:	xpb = 256'h00005800000000000000000000000000000057ffffffa8000000000000005800;
		6'b001100:	xpb = 256'h0000600000000000000000000000000000005fffffffa0000000000000006000;
		6'b001101:	xpb = 256'h00006800000000000000000000000000000067ffffff98000000000000006800;
		6'b001110:	xpb = 256'h0000700000000000000000000000000000006fffffff90000000000000007000;
		6'b001111:	xpb = 256'h00007800000000000000000000000000000077ffffff88000000000000007800;
		6'b010000:	xpb = 256'h0000800000000000000000000000000000007fffffff80000000000000008000;
		6'b010001:	xpb = 256'h00008800000000000000000000000000000087ffffff78000000000000008800;
		6'b010010:	xpb = 256'h0000900000000000000000000000000000008fffffff70000000000000009000;
		6'b010011:	xpb = 256'h00009800000000000000000000000000000097ffffff68000000000000009800;
		6'b010100:	xpb = 256'h0000a00000000000000000000000000000009fffffff6000000000000000a000;
		6'b010101:	xpb = 256'h0000a8000000000000000000000000000000a7ffffff5800000000000000a800;
		6'b010110:	xpb = 256'h0000b0000000000000000000000000000000afffffff5000000000000000b000;
		6'b010111:	xpb = 256'h0000b8000000000000000000000000000000b7ffffff4800000000000000b800;
		6'b011000:	xpb = 256'h0000c0000000000000000000000000000000bfffffff4000000000000000c000;
		6'b011001:	xpb = 256'h0000c8000000000000000000000000000000c7ffffff3800000000000000c800;
		6'b011010:	xpb = 256'h0000d0000000000000000000000000000000cfffffff3000000000000000d000;
		6'b011011:	xpb = 256'h0000d8000000000000000000000000000000d7ffffff2800000000000000d800;
		6'b011100:	xpb = 256'h0000e0000000000000000000000000000000dfffffff2000000000000000e000;
		6'b011101:	xpb = 256'h0000e8000000000000000000000000000000e7ffffff1800000000000000e800;
		6'b011110:	xpb = 256'h0000f0000000000000000000000000000000efffffff1000000000000000f000;
		6'b011111:	xpb = 256'h0000f8000000000000000000000000000000f7ffffff0800000000000000f800;
		6'b100000:	xpb = 256'h000100000000000000000000000000000000ffffffff00000000000000010000;
		6'b100001:	xpb = 256'h00010800000000000000000000000000000107fffffef8000000000000010800;
		6'b100010:	xpb = 256'h0001100000000000000000000000000000010ffffffef0000000000000011000;
		6'b100011:	xpb = 256'h00011800000000000000000000000000000117fffffee8000000000000011800;
		6'b100100:	xpb = 256'h0001200000000000000000000000000000011ffffffee0000000000000012000;
		6'b100101:	xpb = 256'h00012800000000000000000000000000000127fffffed8000000000000012800;
		6'b100110:	xpb = 256'h0001300000000000000000000000000000012ffffffed0000000000000013000;
		6'b100111:	xpb = 256'h00013800000000000000000000000000000137fffffec8000000000000013800;
		6'b101000:	xpb = 256'h0001400000000000000000000000000000013ffffffec0000000000000014000;
		6'b101001:	xpb = 256'h00014800000000000000000000000000000147fffffeb8000000000000014800;
		6'b101010:	xpb = 256'h0001500000000000000000000000000000014ffffffeb0000000000000015000;
		6'b101011:	xpb = 256'h00015800000000000000000000000000000157fffffea8000000000000015800;
		6'b101100:	xpb = 256'h0001600000000000000000000000000000015ffffffea0000000000000016000;
		6'b101101:	xpb = 256'h00016800000000000000000000000000000167fffffe98000000000000016800;
		6'b101110:	xpb = 256'h0001700000000000000000000000000000016ffffffe90000000000000017000;
		6'b101111:	xpb = 256'h00017800000000000000000000000000000177fffffe88000000000000017800;
		6'b110000:	xpb = 256'h0001800000000000000000000000000000017ffffffe80000000000000018000;
		6'b110001:	xpb = 256'h00018800000000000000000000000000000187fffffe78000000000000018800;
		6'b110010:	xpb = 256'h0001900000000000000000000000000000018ffffffe70000000000000019000;
		6'b110011:	xpb = 256'h00019800000000000000000000000000000197fffffe68000000000000019800;
		6'b110100:	xpb = 256'h0001a00000000000000000000000000000019ffffffe6000000000000001a000;
		6'b110101:	xpb = 256'h0001a8000000000000000000000000000001a7fffffe5800000000000001a800;
		6'b110110:	xpb = 256'h0001b0000000000000000000000000000001affffffe5000000000000001b000;
		6'b110111:	xpb = 256'h0001b8000000000000000000000000000001b7fffffe4800000000000001b800;
		6'b111000:	xpb = 256'h0001c0000000000000000000000000000001bffffffe4000000000000001c000;
		6'b111001:	xpb = 256'h0001c8000000000000000000000000000001c7fffffe3800000000000001c800;
		6'b111010:	xpb = 256'h0001d0000000000000000000000000000001cffffffe3000000000000001d000;
		6'b111011:	xpb = 256'h0001d8000000000000000000000000000001d7fffffe2800000000000001d800;
		6'b111100:	xpb = 256'h0001e0000000000000000000000000000001dffffffe2000000000000001e000;
		6'b111101:	xpb = 256'h0001e8000000000000000000000000000001e7fffffe1800000000000001e800;
		6'b111110:	xpb = 256'h0001f0000000000000000000000000000001effffffe1000000000000001f000;
		6'b111111:	xpb = 256'h0001f8000000000000000000000000000001f7fffffe0800000000000001f800;
	endcase
end
endmodule

module xpb_17_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h000100000000000000000000000000000000ffffffff00000000000000010000;
		5'b00010:	xpb = 256'h000200000000000000000000000000000001fffffffe00000000000000020000;
		5'b00011:	xpb = 256'h000300000000000000000000000000000002fffffffd00000000000000030000;
		5'b00100:	xpb = 256'h000400000000000000000000000000000003fffffffc00000000000000040000;
		5'b00101:	xpb = 256'h000500000000000000000000000000000004fffffffb00000000000000050000;
		5'b00110:	xpb = 256'h000600000000000000000000000000000005fffffffa00000000000000060000;
		5'b00111:	xpb = 256'h000700000000000000000000000000000006fffffff900000000000000070000;
		5'b01000:	xpb = 256'h000800000000000000000000000000000007fffffff800000000000000080000;
		5'b01001:	xpb = 256'h000900000000000000000000000000000008fffffff700000000000000090000;
		5'b01010:	xpb = 256'h000a00000000000000000000000000000009fffffff6000000000000000a0000;
		5'b01011:	xpb = 256'h000b0000000000000000000000000000000afffffff5000000000000000b0000;
		5'b01100:	xpb = 256'h000c0000000000000000000000000000000bfffffff4000000000000000c0000;
		5'b01101:	xpb = 256'h000d0000000000000000000000000000000cfffffff3000000000000000d0000;
		5'b01110:	xpb = 256'h000e0000000000000000000000000000000dfffffff2000000000000000e0000;
		5'b01111:	xpb = 256'h000f0000000000000000000000000000000efffffff1000000000000000f0000;
		5'b10000:	xpb = 256'h00100000000000000000000000000000000ffffffff000000000000000100000;
		5'b10001:	xpb = 256'h001100000000000000000000000000000010ffffffef00000000000000110000;
		5'b10010:	xpb = 256'h001200000000000000000000000000000011ffffffee00000000000000120000;
		5'b10011:	xpb = 256'h001300000000000000000000000000000012ffffffed00000000000000130000;
		5'b10100:	xpb = 256'h001400000000000000000000000000000013ffffffec00000000000000140000;
		5'b10101:	xpb = 256'h001500000000000000000000000000000014ffffffeb00000000000000150000;
		5'b10110:	xpb = 256'h001600000000000000000000000000000015ffffffea00000000000000160000;
		5'b10111:	xpb = 256'h001700000000000000000000000000000016ffffffe900000000000000170000;
		5'b11000:	xpb = 256'h001800000000000000000000000000000017ffffffe800000000000000180000;
		5'b11001:	xpb = 256'h001900000000000000000000000000000018ffffffe700000000000000190000;
		5'b11010:	xpb = 256'h001a00000000000000000000000000000019ffffffe6000000000000001a0000;
		5'b11011:	xpb = 256'h001b0000000000000000000000000000001affffffe5000000000000001b0000;
		5'b11100:	xpb = 256'h001c0000000000000000000000000000001bffffffe4000000000000001c0000;
		5'b11101:	xpb = 256'h001d0000000000000000000000000000001cffffffe3000000000000001d0000;
		5'b11110:	xpb = 256'h001e0000000000000000000000000000001dffffffe2000000000000001e0000;
		5'b11111:	xpb = 256'h001f0000000000000000000000000000001effffffe1000000000000001f0000;
	endcase
end
endmodule

module xpb_17_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00200000000000000000000000000000001fffffffe000000000000000200000;
		6'b000010:	xpb = 256'h00400000000000000000000000000000003fffffffc000000000000000400000;
		6'b000011:	xpb = 256'h00600000000000000000000000000000005fffffffa000000000000000600000;
		6'b000100:	xpb = 256'h00800000000000000000000000000000007fffffff8000000000000000800000;
		6'b000101:	xpb = 256'h00a00000000000000000000000000000009fffffff6000000000000000a00000;
		6'b000110:	xpb = 256'h00c0000000000000000000000000000000bfffffff4000000000000000c00000;
		6'b000111:	xpb = 256'h00e0000000000000000000000000000000dfffffff2000000000000000e00000;
		6'b001000:	xpb = 256'h0100000000000000000000000000000000ffffffff0000000000000001000000;
		6'b001001:	xpb = 256'h01200000000000000000000000000000011ffffffee000000000000001200000;
		6'b001010:	xpb = 256'h01400000000000000000000000000000013ffffffec000000000000001400000;
		6'b001011:	xpb = 256'h01600000000000000000000000000000015ffffffea000000000000001600000;
		6'b001100:	xpb = 256'h01800000000000000000000000000000017ffffffe8000000000000001800000;
		6'b001101:	xpb = 256'h01a00000000000000000000000000000019ffffffe6000000000000001a00000;
		6'b001110:	xpb = 256'h01c0000000000000000000000000000001bffffffe4000000000000001c00000;
		6'b001111:	xpb = 256'h01e0000000000000000000000000000001dffffffe2000000000000001e00000;
		6'b010000:	xpb = 256'h0200000000000000000000000000000001fffffffe0000000000000002000000;
		6'b010001:	xpb = 256'h02200000000000000000000000000000021ffffffde000000000000002200000;
		6'b010010:	xpb = 256'h02400000000000000000000000000000023ffffffdc000000000000002400000;
		6'b010011:	xpb = 256'h02600000000000000000000000000000025ffffffda000000000000002600000;
		6'b010100:	xpb = 256'h02800000000000000000000000000000027ffffffd8000000000000002800000;
		6'b010101:	xpb = 256'h02a00000000000000000000000000000029ffffffd6000000000000002a00000;
		6'b010110:	xpb = 256'h02c0000000000000000000000000000002bffffffd4000000000000002c00000;
		6'b010111:	xpb = 256'h02e0000000000000000000000000000002dffffffd2000000000000002e00000;
		6'b011000:	xpb = 256'h0300000000000000000000000000000002fffffffd0000000000000003000000;
		6'b011001:	xpb = 256'h03200000000000000000000000000000031ffffffce000000000000003200000;
		6'b011010:	xpb = 256'h03400000000000000000000000000000033ffffffcc000000000000003400000;
		6'b011011:	xpb = 256'h03600000000000000000000000000000035ffffffca000000000000003600000;
		6'b011100:	xpb = 256'h03800000000000000000000000000000037ffffffc8000000000000003800000;
		6'b011101:	xpb = 256'h03a00000000000000000000000000000039ffffffc6000000000000003a00000;
		6'b011110:	xpb = 256'h03c0000000000000000000000000000003bffffffc4000000000000003c00000;
		6'b011111:	xpb = 256'h03e0000000000000000000000000000003dffffffc2000000000000003e00000;
		6'b100000:	xpb = 256'h0400000000000000000000000000000003fffffffc0000000000000004000000;
		6'b100001:	xpb = 256'h04200000000000000000000000000000041ffffffbe000000000000004200000;
		6'b100010:	xpb = 256'h04400000000000000000000000000000043ffffffbc000000000000004400000;
		6'b100011:	xpb = 256'h04600000000000000000000000000000045ffffffba000000000000004600000;
		6'b100100:	xpb = 256'h04800000000000000000000000000000047ffffffb8000000000000004800000;
		6'b100101:	xpb = 256'h04a00000000000000000000000000000049ffffffb6000000000000004a00000;
		6'b100110:	xpb = 256'h04c0000000000000000000000000000004bffffffb4000000000000004c00000;
		6'b100111:	xpb = 256'h04e0000000000000000000000000000004dffffffb2000000000000004e00000;
		6'b101000:	xpb = 256'h0500000000000000000000000000000004fffffffb0000000000000005000000;
		6'b101001:	xpb = 256'h05200000000000000000000000000000051ffffffae000000000000005200000;
		6'b101010:	xpb = 256'h05400000000000000000000000000000053ffffffac000000000000005400000;
		6'b101011:	xpb = 256'h05600000000000000000000000000000055ffffffaa000000000000005600000;
		6'b101100:	xpb = 256'h05800000000000000000000000000000057ffffffa8000000000000005800000;
		6'b101101:	xpb = 256'h05a00000000000000000000000000000059ffffffa6000000000000005a00000;
		6'b101110:	xpb = 256'h05c0000000000000000000000000000005bffffffa4000000000000005c00000;
		6'b101111:	xpb = 256'h05e0000000000000000000000000000005dffffffa2000000000000005e00000;
		6'b110000:	xpb = 256'h0600000000000000000000000000000005fffffffa0000000000000006000000;
		6'b110001:	xpb = 256'h06200000000000000000000000000000061ffffff9e000000000000006200000;
		6'b110010:	xpb = 256'h06400000000000000000000000000000063ffffff9c000000000000006400000;
		6'b110011:	xpb = 256'h06600000000000000000000000000000065ffffff9a000000000000006600000;
		6'b110100:	xpb = 256'h06800000000000000000000000000000067ffffff98000000000000006800000;
		6'b110101:	xpb = 256'h06a00000000000000000000000000000069ffffff96000000000000006a00000;
		6'b110110:	xpb = 256'h06c0000000000000000000000000000006bffffff94000000000000006c00000;
		6'b110111:	xpb = 256'h06e0000000000000000000000000000006dffffff92000000000000006e00000;
		6'b111000:	xpb = 256'h0700000000000000000000000000000006fffffff90000000000000007000000;
		6'b111001:	xpb = 256'h07200000000000000000000000000000071ffffff8e000000000000007200000;
		6'b111010:	xpb = 256'h07400000000000000000000000000000073ffffff8c000000000000007400000;
		6'b111011:	xpb = 256'h07600000000000000000000000000000075ffffff8a000000000000007600000;
		6'b111100:	xpb = 256'h07800000000000000000000000000000077ffffff88000000000000007800000;
		6'b111101:	xpb = 256'h07a00000000000000000000000000000079ffffff86000000000000007a00000;
		6'b111110:	xpb = 256'h07c0000000000000000000000000000007bffffff84000000000000007c00000;
		6'b111111:	xpb = 256'h07e0000000000000000000000000000007dffffff82000000000000007e00000;
	endcase
end
endmodule

module xpb_17_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0800000000000000000000000000000007fffffff80000000000000008000000;
		6'b000010:	xpb = 256'h100000000000000000000000000000000ffffffff00000000000000010000000;
		6'b000011:	xpb = 256'h1800000000000000000000000000000017ffffffe80000000000000018000000;
		6'b000100:	xpb = 256'h200000000000000000000000000000001fffffffe00000000000000020000000;
		6'b000101:	xpb = 256'h2800000000000000000000000000000027ffffffd80000000000000028000000;
		6'b000110:	xpb = 256'h300000000000000000000000000000002fffffffd00000000000000030000000;
		6'b000111:	xpb = 256'h3800000000000000000000000000000037ffffffc80000000000000038000000;
		6'b001000:	xpb = 256'h400000000000000000000000000000003fffffffc00000000000000040000000;
		6'b001001:	xpb = 256'h4800000000000000000000000000000047ffffffb80000000000000048000000;
		6'b001010:	xpb = 256'h500000000000000000000000000000004fffffffb00000000000000050000000;
		6'b001011:	xpb = 256'h5800000000000000000000000000000057ffffffa80000000000000058000000;
		6'b001100:	xpb = 256'h600000000000000000000000000000005fffffffa00000000000000060000000;
		6'b001101:	xpb = 256'h6800000000000000000000000000000067ffffff980000000000000068000000;
		6'b001110:	xpb = 256'h700000000000000000000000000000006fffffff900000000000000070000000;
		6'b001111:	xpb = 256'h7800000000000000000000000000000077ffffff880000000000000078000000;
		6'b010000:	xpb = 256'h800000000000000000000000000000007fffffff800000000000000080000000;
		6'b010001:	xpb = 256'h8800000000000000000000000000000087ffffff780000000000000088000000;
		6'b010010:	xpb = 256'h900000000000000000000000000000008fffffff700000000000000090000000;
		6'b010011:	xpb = 256'h9800000000000000000000000000000097ffffff680000000000000098000000;
		6'b010100:	xpb = 256'ha00000000000000000000000000000009fffffff6000000000000000a0000000;
		6'b010101:	xpb = 256'ha8000000000000000000000000000000a7ffffff5800000000000000a8000000;
		6'b010110:	xpb = 256'hb0000000000000000000000000000000afffffff5000000000000000b0000000;
		6'b010111:	xpb = 256'hb8000000000000000000000000000000b7ffffff4800000000000000b8000000;
		6'b011000:	xpb = 256'hc0000000000000000000000000000000bfffffff4000000000000000c0000000;
		6'b011001:	xpb = 256'hc8000000000000000000000000000000c7ffffff3800000000000000c8000000;
		6'b011010:	xpb = 256'hd0000000000000000000000000000000cfffffff3000000000000000d0000000;
		6'b011011:	xpb = 256'hd8000000000000000000000000000000d7ffffff2800000000000000d8000000;
		6'b011100:	xpb = 256'he0000000000000000000000000000000dfffffff2000000000000000e0000000;
		6'b011101:	xpb = 256'he8000000000000000000000000000000e7ffffff1800000000000000e8000000;
		6'b011110:	xpb = 256'hf0000000000000000000000000000000efffffff1000000000000000f0000000;
		6'b011111:	xpb = 256'hf8000000000000000000000000000000f7ffffff0800000000000000f8000000;
		6'b100000:	xpb = 256'h00000001000000000000000000000000ffffffffffffffff0000000100000001;
		6'b100001:	xpb = 256'h0800000100000000000000000000000107fffffff7ffffff0000000108000001;
		6'b100010:	xpb = 256'h100000010000000000000000000000010fffffffefffffff0000000110000001;
		6'b100011:	xpb = 256'h1800000100000000000000000000000117ffffffe7ffffff0000000118000001;
		6'b100100:	xpb = 256'h200000010000000000000000000000011fffffffdfffffff0000000120000001;
		6'b100101:	xpb = 256'h2800000100000000000000000000000127ffffffd7ffffff0000000128000001;
		6'b100110:	xpb = 256'h300000010000000000000000000000012fffffffcfffffff0000000130000001;
		6'b100111:	xpb = 256'h3800000100000000000000000000000137ffffffc7ffffff0000000138000001;
		6'b101000:	xpb = 256'h400000010000000000000000000000013fffffffbfffffff0000000140000001;
		6'b101001:	xpb = 256'h4800000100000000000000000000000147ffffffb7ffffff0000000148000001;
		6'b101010:	xpb = 256'h500000010000000000000000000000014fffffffafffffff0000000150000001;
		6'b101011:	xpb = 256'h5800000100000000000000000000000157ffffffa7ffffff0000000158000001;
		6'b101100:	xpb = 256'h600000010000000000000000000000015fffffff9fffffff0000000160000001;
		6'b101101:	xpb = 256'h6800000100000000000000000000000167ffffff97ffffff0000000168000001;
		6'b101110:	xpb = 256'h700000010000000000000000000000016fffffff8fffffff0000000170000001;
		6'b101111:	xpb = 256'h7800000100000000000000000000000177ffffff87ffffff0000000178000001;
		6'b110000:	xpb = 256'h800000010000000000000000000000017fffffff7fffffff0000000180000001;
		6'b110001:	xpb = 256'h8800000100000000000000000000000187ffffff77ffffff0000000188000001;
		6'b110010:	xpb = 256'h900000010000000000000000000000018fffffff6fffffff0000000190000001;
		6'b110011:	xpb = 256'h9800000100000000000000000000000197ffffff67ffffff0000000198000001;
		6'b110100:	xpb = 256'ha00000010000000000000000000000019fffffff5fffffff00000001a0000001;
		6'b110101:	xpb = 256'ha8000001000000000000000000000001a7ffffff57ffffff00000001a8000001;
		6'b110110:	xpb = 256'hb0000001000000000000000000000001afffffff4fffffff00000001b0000001;
		6'b110111:	xpb = 256'hb8000001000000000000000000000001b7ffffff47ffffff00000001b8000001;
		6'b111000:	xpb = 256'hc0000001000000000000000000000001bfffffff3fffffff00000001c0000001;
		6'b111001:	xpb = 256'hc8000001000000000000000000000001c7ffffff37ffffff00000001c8000001;
		6'b111010:	xpb = 256'hd0000001000000000000000000000001cfffffff2fffffff00000001d0000001;
		6'b111011:	xpb = 256'hd8000001000000000000000000000001d7ffffff27ffffff00000001d8000001;
		6'b111100:	xpb = 256'he0000001000000000000000000000001dfffffff1fffffff00000001e0000001;
		6'b111101:	xpb = 256'he8000001000000000000000000000001e7ffffff17ffffff00000001e8000001;
		6'b111110:	xpb = 256'hf0000001000000000000000000000001efffffff0fffffff00000001f0000001;
		6'b111111:	xpb = 256'hf8000001000000000000000000000001f7ffffff07ffffff00000001f8000001;
	endcase
end
endmodule

module xpb_18_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h00000001000000000000000000000000ffffffffffffffff0000000100000001;
		5'b00010:	xpb = 256'h00000002000000000000000000000001fffffffffffffffe0000000200000002;
		5'b00011:	xpb = 256'h00000003000000000000000000000002fffffffffffffffd0000000300000003;
		5'b00100:	xpb = 256'h00000004000000000000000000000003fffffffffffffffc0000000400000004;
		5'b00101:	xpb = 256'h00000005000000000000000000000004fffffffffffffffb0000000500000005;
		5'b00110:	xpb = 256'h00000006000000000000000000000005fffffffffffffffa0000000600000006;
		5'b00111:	xpb = 256'h00000007000000000000000000000006fffffffffffffff90000000700000007;
		5'b01000:	xpb = 256'h00000008000000000000000000000007fffffffffffffff80000000800000008;
		5'b01001:	xpb = 256'h00000009000000000000000000000008fffffffffffffff70000000900000009;
		5'b01010:	xpb = 256'h0000000a000000000000000000000009fffffffffffffff60000000a0000000a;
		5'b01011:	xpb = 256'h0000000b00000000000000000000000afffffffffffffff50000000b0000000b;
		5'b01100:	xpb = 256'h0000000c00000000000000000000000bfffffffffffffff40000000c0000000c;
		5'b01101:	xpb = 256'h0000000d00000000000000000000000cfffffffffffffff30000000d0000000d;
		5'b01110:	xpb = 256'h0000000e00000000000000000000000dfffffffffffffff20000000e0000000e;
		5'b01111:	xpb = 256'h0000000f00000000000000000000000efffffffffffffff10000000f0000000f;
		5'b10000:	xpb = 256'h0000001000000000000000000000000ffffffffffffffff00000001000000010;
		5'b10001:	xpb = 256'h00000011000000000000000000000010ffffffffffffffef0000001100000011;
		5'b10010:	xpb = 256'h00000012000000000000000000000011ffffffffffffffee0000001200000012;
		5'b10011:	xpb = 256'h00000013000000000000000000000012ffffffffffffffed0000001300000013;
		5'b10100:	xpb = 256'h00000014000000000000000000000013ffffffffffffffec0000001400000014;
		5'b10101:	xpb = 256'h00000015000000000000000000000014ffffffffffffffeb0000001500000015;
		5'b10110:	xpb = 256'h00000016000000000000000000000015ffffffffffffffea0000001600000016;
		5'b10111:	xpb = 256'h00000017000000000000000000000016ffffffffffffffe90000001700000017;
		5'b11000:	xpb = 256'h00000018000000000000000000000017ffffffffffffffe80000001800000018;
		5'b11001:	xpb = 256'h00000019000000000000000000000018ffffffffffffffe70000001900000019;
		5'b11010:	xpb = 256'h0000001a000000000000000000000019ffffffffffffffe60000001a0000001a;
		5'b11011:	xpb = 256'h0000001b00000000000000000000001affffffffffffffe50000001b0000001b;
		5'b11100:	xpb = 256'h0000001c00000000000000000000001bffffffffffffffe40000001c0000001c;
		5'b11101:	xpb = 256'h0000001d00000000000000000000001cffffffffffffffe30000001d0000001d;
		5'b11110:	xpb = 256'h0000001e00000000000000000000001dffffffffffffffe20000001e0000001e;
		5'b11111:	xpb = 256'h0000001f00000000000000000000001effffffffffffffe10000001f0000001f;
	endcase
end
endmodule

module xpb_18_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000002000000000000000000000001fffffffffffffffe00000002000000020;
		6'b000010:	xpb = 256'h0000004000000000000000000000003fffffffffffffffc00000004000000040;
		6'b000011:	xpb = 256'h0000006000000000000000000000005fffffffffffffffa00000006000000060;
		6'b000100:	xpb = 256'h0000008000000000000000000000007fffffffffffffff800000008000000080;
		6'b000101:	xpb = 256'h000000a000000000000000000000009fffffffffffffff60000000a0000000a0;
		6'b000110:	xpb = 256'h000000c00000000000000000000000bfffffffffffffff40000000c0000000c0;
		6'b000111:	xpb = 256'h000000e00000000000000000000000dfffffffffffffff20000000e0000000e0;
		6'b001000:	xpb = 256'h000001000000000000000000000000ffffffffffffffff000000010000000100;
		6'b001001:	xpb = 256'h0000012000000000000000000000011ffffffffffffffee00000012000000120;
		6'b001010:	xpb = 256'h0000014000000000000000000000013ffffffffffffffec00000014000000140;
		6'b001011:	xpb = 256'h0000016000000000000000000000015ffffffffffffffea00000016000000160;
		6'b001100:	xpb = 256'h0000018000000000000000000000017ffffffffffffffe800000018000000180;
		6'b001101:	xpb = 256'h000001a000000000000000000000019ffffffffffffffe60000001a0000001a0;
		6'b001110:	xpb = 256'h000001c00000000000000000000001bffffffffffffffe40000001c0000001c0;
		6'b001111:	xpb = 256'h000001e00000000000000000000001dffffffffffffffe20000001e0000001e0;
		6'b010000:	xpb = 256'h000002000000000000000000000001fffffffffffffffe000000020000000200;
		6'b010001:	xpb = 256'h0000022000000000000000000000021ffffffffffffffde00000022000000220;
		6'b010010:	xpb = 256'h0000024000000000000000000000023ffffffffffffffdc00000024000000240;
		6'b010011:	xpb = 256'h0000026000000000000000000000025ffffffffffffffda00000026000000260;
		6'b010100:	xpb = 256'h0000028000000000000000000000027ffffffffffffffd800000028000000280;
		6'b010101:	xpb = 256'h000002a000000000000000000000029ffffffffffffffd60000002a0000002a0;
		6'b010110:	xpb = 256'h000002c00000000000000000000002bffffffffffffffd40000002c0000002c0;
		6'b010111:	xpb = 256'h000002e00000000000000000000002dffffffffffffffd20000002e0000002e0;
		6'b011000:	xpb = 256'h000003000000000000000000000002fffffffffffffffd000000030000000300;
		6'b011001:	xpb = 256'h0000032000000000000000000000031ffffffffffffffce00000032000000320;
		6'b011010:	xpb = 256'h0000034000000000000000000000033ffffffffffffffcc00000034000000340;
		6'b011011:	xpb = 256'h0000036000000000000000000000035ffffffffffffffca00000036000000360;
		6'b011100:	xpb = 256'h0000038000000000000000000000037ffffffffffffffc800000038000000380;
		6'b011101:	xpb = 256'h000003a000000000000000000000039ffffffffffffffc60000003a0000003a0;
		6'b011110:	xpb = 256'h000003c00000000000000000000003bffffffffffffffc40000003c0000003c0;
		6'b011111:	xpb = 256'h000003e00000000000000000000003dffffffffffffffc20000003e0000003e0;
		6'b100000:	xpb = 256'h000004000000000000000000000003fffffffffffffffc000000040000000400;
		6'b100001:	xpb = 256'h0000042000000000000000000000041ffffffffffffffbe00000042000000420;
		6'b100010:	xpb = 256'h0000044000000000000000000000043ffffffffffffffbc00000044000000440;
		6'b100011:	xpb = 256'h0000046000000000000000000000045ffffffffffffffba00000046000000460;
		6'b100100:	xpb = 256'h0000048000000000000000000000047ffffffffffffffb800000048000000480;
		6'b100101:	xpb = 256'h000004a000000000000000000000049ffffffffffffffb60000004a0000004a0;
		6'b100110:	xpb = 256'h000004c00000000000000000000004bffffffffffffffb40000004c0000004c0;
		6'b100111:	xpb = 256'h000004e00000000000000000000004dffffffffffffffb20000004e0000004e0;
		6'b101000:	xpb = 256'h000005000000000000000000000004fffffffffffffffb000000050000000500;
		6'b101001:	xpb = 256'h0000052000000000000000000000051ffffffffffffffae00000052000000520;
		6'b101010:	xpb = 256'h0000054000000000000000000000053ffffffffffffffac00000054000000540;
		6'b101011:	xpb = 256'h0000056000000000000000000000055ffffffffffffffaa00000056000000560;
		6'b101100:	xpb = 256'h0000058000000000000000000000057ffffffffffffffa800000058000000580;
		6'b101101:	xpb = 256'h000005a000000000000000000000059ffffffffffffffa60000005a0000005a0;
		6'b101110:	xpb = 256'h000005c00000000000000000000005bffffffffffffffa40000005c0000005c0;
		6'b101111:	xpb = 256'h000005e00000000000000000000005dffffffffffffffa20000005e0000005e0;
		6'b110000:	xpb = 256'h000006000000000000000000000005fffffffffffffffa000000060000000600;
		6'b110001:	xpb = 256'h0000062000000000000000000000061ffffffffffffff9e00000062000000620;
		6'b110010:	xpb = 256'h0000064000000000000000000000063ffffffffffffff9c00000064000000640;
		6'b110011:	xpb = 256'h0000066000000000000000000000065ffffffffffffff9a00000066000000660;
		6'b110100:	xpb = 256'h0000068000000000000000000000067ffffffffffffff9800000068000000680;
		6'b110101:	xpb = 256'h000006a000000000000000000000069ffffffffffffff960000006a0000006a0;
		6'b110110:	xpb = 256'h000006c00000000000000000000006bffffffffffffff940000006c0000006c0;
		6'b110111:	xpb = 256'h000006e00000000000000000000006dffffffffffffff920000006e0000006e0;
		6'b111000:	xpb = 256'h000007000000000000000000000006fffffffffffffff9000000070000000700;
		6'b111001:	xpb = 256'h0000072000000000000000000000071ffffffffffffff8e00000072000000720;
		6'b111010:	xpb = 256'h0000074000000000000000000000073ffffffffffffff8c00000074000000740;
		6'b111011:	xpb = 256'h0000076000000000000000000000075ffffffffffffff8a00000076000000760;
		6'b111100:	xpb = 256'h0000078000000000000000000000077ffffffffffffff8800000078000000780;
		6'b111101:	xpb = 256'h000007a000000000000000000000079ffffffffffffff860000007a0000007a0;
		6'b111110:	xpb = 256'h000007c00000000000000000000007bffffffffffffff840000007c0000007c0;
		6'b111111:	xpb = 256'h000007e00000000000000000000007dffffffffffffff820000007e0000007e0;
	endcase
end
endmodule

module xpb_18_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h000008000000000000000000000007fffffffffffffff8000000080000000800;
		6'b000010:	xpb = 256'h00001000000000000000000000000ffffffffffffffff0000000100000001000;
		6'b000011:	xpb = 256'h000018000000000000000000000017ffffffffffffffe8000000180000001800;
		6'b000100:	xpb = 256'h00002000000000000000000000001fffffffffffffffe0000000200000002000;
		6'b000101:	xpb = 256'h000028000000000000000000000027ffffffffffffffd8000000280000002800;
		6'b000110:	xpb = 256'h00003000000000000000000000002fffffffffffffffd0000000300000003000;
		6'b000111:	xpb = 256'h000038000000000000000000000037ffffffffffffffc8000000380000003800;
		6'b001000:	xpb = 256'h00004000000000000000000000003fffffffffffffffc0000000400000004000;
		6'b001001:	xpb = 256'h000048000000000000000000000047ffffffffffffffb8000000480000004800;
		6'b001010:	xpb = 256'h00005000000000000000000000004fffffffffffffffb0000000500000005000;
		6'b001011:	xpb = 256'h000058000000000000000000000057ffffffffffffffa8000000580000005800;
		6'b001100:	xpb = 256'h00006000000000000000000000005fffffffffffffffa0000000600000006000;
		6'b001101:	xpb = 256'h000068000000000000000000000067ffffffffffffff98000000680000006800;
		6'b001110:	xpb = 256'h00007000000000000000000000006fffffffffffffff90000000700000007000;
		6'b001111:	xpb = 256'h000078000000000000000000000077ffffffffffffff88000000780000007800;
		6'b010000:	xpb = 256'h00008000000000000000000000007fffffffffffffff80000000800000008000;
		6'b010001:	xpb = 256'h000088000000000000000000000087ffffffffffffff78000000880000008800;
		6'b010010:	xpb = 256'h00009000000000000000000000008fffffffffffffff70000000900000009000;
		6'b010011:	xpb = 256'h000098000000000000000000000097ffffffffffffff68000000980000009800;
		6'b010100:	xpb = 256'h0000a000000000000000000000009fffffffffffffff60000000a0000000a000;
		6'b010101:	xpb = 256'h0000a80000000000000000000000a7ffffffffffffff58000000a8000000a800;
		6'b010110:	xpb = 256'h0000b00000000000000000000000afffffffffffffff50000000b0000000b000;
		6'b010111:	xpb = 256'h0000b80000000000000000000000b7ffffffffffffff48000000b8000000b800;
		6'b011000:	xpb = 256'h0000c00000000000000000000000bfffffffffffffff40000000c0000000c000;
		6'b011001:	xpb = 256'h0000c80000000000000000000000c7ffffffffffffff38000000c8000000c800;
		6'b011010:	xpb = 256'h0000d00000000000000000000000cfffffffffffffff30000000d0000000d000;
		6'b011011:	xpb = 256'h0000d80000000000000000000000d7ffffffffffffff28000000d8000000d800;
		6'b011100:	xpb = 256'h0000e00000000000000000000000dfffffffffffffff20000000e0000000e000;
		6'b011101:	xpb = 256'h0000e80000000000000000000000e7ffffffffffffff18000000e8000000e800;
		6'b011110:	xpb = 256'h0000f00000000000000000000000efffffffffffffff10000000f0000000f000;
		6'b011111:	xpb = 256'h0000f80000000000000000000000f7ffffffffffffff08000000f8000000f800;
		6'b100000:	xpb = 256'h0001000000000000000000000000ffffffffffffffff00000001000000010000;
		6'b100001:	xpb = 256'h000108000000000000000000000107fffffffffffffef8000001080000010800;
		6'b100010:	xpb = 256'h00011000000000000000000000010ffffffffffffffef0000001100000011000;
		6'b100011:	xpb = 256'h000118000000000000000000000117fffffffffffffee8000001180000011800;
		6'b100100:	xpb = 256'h00012000000000000000000000011ffffffffffffffee0000001200000012000;
		6'b100101:	xpb = 256'h000128000000000000000000000127fffffffffffffed8000001280000012800;
		6'b100110:	xpb = 256'h00013000000000000000000000012ffffffffffffffed0000001300000013000;
		6'b100111:	xpb = 256'h000138000000000000000000000137fffffffffffffec8000001380000013800;
		6'b101000:	xpb = 256'h00014000000000000000000000013ffffffffffffffec0000001400000014000;
		6'b101001:	xpb = 256'h000148000000000000000000000147fffffffffffffeb8000001480000014800;
		6'b101010:	xpb = 256'h00015000000000000000000000014ffffffffffffffeb0000001500000015000;
		6'b101011:	xpb = 256'h000158000000000000000000000157fffffffffffffea8000001580000015800;
		6'b101100:	xpb = 256'h00016000000000000000000000015ffffffffffffffea0000001600000016000;
		6'b101101:	xpb = 256'h000168000000000000000000000167fffffffffffffe98000001680000016800;
		6'b101110:	xpb = 256'h00017000000000000000000000016ffffffffffffffe90000001700000017000;
		6'b101111:	xpb = 256'h000178000000000000000000000177fffffffffffffe88000001780000017800;
		6'b110000:	xpb = 256'h00018000000000000000000000017ffffffffffffffe80000001800000018000;
		6'b110001:	xpb = 256'h000188000000000000000000000187fffffffffffffe78000001880000018800;
		6'b110010:	xpb = 256'h00019000000000000000000000018ffffffffffffffe70000001900000019000;
		6'b110011:	xpb = 256'h000198000000000000000000000197fffffffffffffe68000001980000019800;
		6'b110100:	xpb = 256'h0001a000000000000000000000019ffffffffffffffe60000001a0000001a000;
		6'b110101:	xpb = 256'h0001a80000000000000000000001a7fffffffffffffe58000001a8000001a800;
		6'b110110:	xpb = 256'h0001b00000000000000000000001affffffffffffffe50000001b0000001b000;
		6'b110111:	xpb = 256'h0001b80000000000000000000001b7fffffffffffffe48000001b8000001b800;
		6'b111000:	xpb = 256'h0001c00000000000000000000001bffffffffffffffe40000001c0000001c000;
		6'b111001:	xpb = 256'h0001c80000000000000000000001c7fffffffffffffe38000001c8000001c800;
		6'b111010:	xpb = 256'h0001d00000000000000000000001cffffffffffffffe30000001d0000001d000;
		6'b111011:	xpb = 256'h0001d80000000000000000000001d7fffffffffffffe28000001d8000001d800;
		6'b111100:	xpb = 256'h0001e00000000000000000000001dffffffffffffffe20000001e0000001e000;
		6'b111101:	xpb = 256'h0001e80000000000000000000001e7fffffffffffffe18000001e8000001e800;
		6'b111110:	xpb = 256'h0001f00000000000000000000001effffffffffffffe10000001f0000001f000;
		6'b111111:	xpb = 256'h0001f80000000000000000000001f7fffffffffffffe08000001f8000001f800;
	endcase
end
endmodule

module xpb_19_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0001000000000000000000000000ffffffffffffffff00000001000000010000;
		5'b00010:	xpb = 256'h0002000000000000000000000001fffffffffffffffe00000002000000020000;
		5'b00011:	xpb = 256'h0003000000000000000000000002fffffffffffffffd00000003000000030000;
		5'b00100:	xpb = 256'h0004000000000000000000000003fffffffffffffffc00000004000000040000;
		5'b00101:	xpb = 256'h0005000000000000000000000004fffffffffffffffb00000005000000050000;
		5'b00110:	xpb = 256'h0006000000000000000000000005fffffffffffffffa00000006000000060000;
		5'b00111:	xpb = 256'h0007000000000000000000000006fffffffffffffff900000007000000070000;
		5'b01000:	xpb = 256'h0008000000000000000000000007fffffffffffffff800000008000000080000;
		5'b01001:	xpb = 256'h0009000000000000000000000008fffffffffffffff700000009000000090000;
		5'b01010:	xpb = 256'h000a000000000000000000000009fffffffffffffff60000000a0000000a0000;
		5'b01011:	xpb = 256'h000b00000000000000000000000afffffffffffffff50000000b0000000b0000;
		5'b01100:	xpb = 256'h000c00000000000000000000000bfffffffffffffff40000000c0000000c0000;
		5'b01101:	xpb = 256'h000d00000000000000000000000cfffffffffffffff30000000d0000000d0000;
		5'b01110:	xpb = 256'h000e00000000000000000000000dfffffffffffffff20000000e0000000e0000;
		5'b01111:	xpb = 256'h000f00000000000000000000000efffffffffffffff10000000f0000000f0000;
		5'b10000:	xpb = 256'h001000000000000000000000000ffffffffffffffff000000010000000100000;
		5'b10001:	xpb = 256'h0011000000000000000000000010ffffffffffffffef00000011000000110000;
		5'b10010:	xpb = 256'h0012000000000000000000000011ffffffffffffffee00000012000000120000;
		5'b10011:	xpb = 256'h0013000000000000000000000012ffffffffffffffed00000013000000130000;
		5'b10100:	xpb = 256'h0014000000000000000000000013ffffffffffffffec00000014000000140000;
		5'b10101:	xpb = 256'h0015000000000000000000000014ffffffffffffffeb00000015000000150000;
		5'b10110:	xpb = 256'h0016000000000000000000000015ffffffffffffffea00000016000000160000;
		5'b10111:	xpb = 256'h0017000000000000000000000016ffffffffffffffe900000017000000170000;
		5'b11000:	xpb = 256'h0018000000000000000000000017ffffffffffffffe800000018000000180000;
		5'b11001:	xpb = 256'h0019000000000000000000000018ffffffffffffffe700000019000000190000;
		5'b11010:	xpb = 256'h001a000000000000000000000019ffffffffffffffe60000001a0000001a0000;
		5'b11011:	xpb = 256'h001b00000000000000000000001affffffffffffffe50000001b0000001b0000;
		5'b11100:	xpb = 256'h001c00000000000000000000001bffffffffffffffe40000001c0000001c0000;
		5'b11101:	xpb = 256'h001d00000000000000000000001cffffffffffffffe30000001d0000001d0000;
		5'b11110:	xpb = 256'h001e00000000000000000000001dffffffffffffffe20000001e0000001e0000;
		5'b11111:	xpb = 256'h001f00000000000000000000001effffffffffffffe10000001f0000001f0000;
	endcase
end
endmodule

module xpb_19_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h002000000000000000000000001fffffffffffffffe000000020000000200000;
		6'b000010:	xpb = 256'h004000000000000000000000003fffffffffffffffc000000040000000400000;
		6'b000011:	xpb = 256'h006000000000000000000000005fffffffffffffffa000000060000000600000;
		6'b000100:	xpb = 256'h008000000000000000000000007fffffffffffffff8000000080000000800000;
		6'b000101:	xpb = 256'h00a000000000000000000000009fffffffffffffff60000000a0000000a00000;
		6'b000110:	xpb = 256'h00c00000000000000000000000bfffffffffffffff40000000c0000000c00000;
		6'b000111:	xpb = 256'h00e00000000000000000000000dfffffffffffffff20000000e0000000e00000;
		6'b001000:	xpb = 256'h01000000000000000000000000ffffffffffffffff0000000100000001000000;
		6'b001001:	xpb = 256'h012000000000000000000000011ffffffffffffffee000000120000001200000;
		6'b001010:	xpb = 256'h014000000000000000000000013ffffffffffffffec000000140000001400000;
		6'b001011:	xpb = 256'h016000000000000000000000015ffffffffffffffea000000160000001600000;
		6'b001100:	xpb = 256'h018000000000000000000000017ffffffffffffffe8000000180000001800000;
		6'b001101:	xpb = 256'h01a000000000000000000000019ffffffffffffffe60000001a0000001a00000;
		6'b001110:	xpb = 256'h01c00000000000000000000001bffffffffffffffe40000001c0000001c00000;
		6'b001111:	xpb = 256'h01e00000000000000000000001dffffffffffffffe20000001e0000001e00000;
		6'b010000:	xpb = 256'h02000000000000000000000001fffffffffffffffe0000000200000002000000;
		6'b010001:	xpb = 256'h022000000000000000000000021ffffffffffffffde000000220000002200000;
		6'b010010:	xpb = 256'h024000000000000000000000023ffffffffffffffdc000000240000002400000;
		6'b010011:	xpb = 256'h026000000000000000000000025ffffffffffffffda000000260000002600000;
		6'b010100:	xpb = 256'h028000000000000000000000027ffffffffffffffd8000000280000002800000;
		6'b010101:	xpb = 256'h02a000000000000000000000029ffffffffffffffd60000002a0000002a00000;
		6'b010110:	xpb = 256'h02c00000000000000000000002bffffffffffffffd40000002c0000002c00000;
		6'b010111:	xpb = 256'h02e00000000000000000000002dffffffffffffffd20000002e0000002e00000;
		6'b011000:	xpb = 256'h03000000000000000000000002fffffffffffffffd0000000300000003000000;
		6'b011001:	xpb = 256'h032000000000000000000000031ffffffffffffffce000000320000003200000;
		6'b011010:	xpb = 256'h034000000000000000000000033ffffffffffffffcc000000340000003400000;
		6'b011011:	xpb = 256'h036000000000000000000000035ffffffffffffffca000000360000003600000;
		6'b011100:	xpb = 256'h038000000000000000000000037ffffffffffffffc8000000380000003800000;
		6'b011101:	xpb = 256'h03a000000000000000000000039ffffffffffffffc60000003a0000003a00000;
		6'b011110:	xpb = 256'h03c00000000000000000000003bffffffffffffffc40000003c0000003c00000;
		6'b011111:	xpb = 256'h03e00000000000000000000003dffffffffffffffc20000003e0000003e00000;
		6'b100000:	xpb = 256'h04000000000000000000000003fffffffffffffffc0000000400000004000000;
		6'b100001:	xpb = 256'h042000000000000000000000041ffffffffffffffbe000000420000004200000;
		6'b100010:	xpb = 256'h044000000000000000000000043ffffffffffffffbc000000440000004400000;
		6'b100011:	xpb = 256'h046000000000000000000000045ffffffffffffffba000000460000004600000;
		6'b100100:	xpb = 256'h048000000000000000000000047ffffffffffffffb8000000480000004800000;
		6'b100101:	xpb = 256'h04a000000000000000000000049ffffffffffffffb60000004a0000004a00000;
		6'b100110:	xpb = 256'h04c00000000000000000000004bffffffffffffffb40000004c0000004c00000;
		6'b100111:	xpb = 256'h04e00000000000000000000004dffffffffffffffb20000004e0000004e00000;
		6'b101000:	xpb = 256'h05000000000000000000000004fffffffffffffffb0000000500000005000000;
		6'b101001:	xpb = 256'h052000000000000000000000051ffffffffffffffae000000520000005200000;
		6'b101010:	xpb = 256'h054000000000000000000000053ffffffffffffffac000000540000005400000;
		6'b101011:	xpb = 256'h056000000000000000000000055ffffffffffffffaa000000560000005600000;
		6'b101100:	xpb = 256'h058000000000000000000000057ffffffffffffffa8000000580000005800000;
		6'b101101:	xpb = 256'h05a000000000000000000000059ffffffffffffffa60000005a0000005a00000;
		6'b101110:	xpb = 256'h05c00000000000000000000005bffffffffffffffa40000005c0000005c00000;
		6'b101111:	xpb = 256'h05e00000000000000000000005dffffffffffffffa20000005e0000005e00000;
		6'b110000:	xpb = 256'h06000000000000000000000005fffffffffffffffa0000000600000006000000;
		6'b110001:	xpb = 256'h062000000000000000000000061ffffffffffffff9e000000620000006200000;
		6'b110010:	xpb = 256'h064000000000000000000000063ffffffffffffff9c000000640000006400000;
		6'b110011:	xpb = 256'h066000000000000000000000065ffffffffffffff9a000000660000006600000;
		6'b110100:	xpb = 256'h068000000000000000000000067ffffffffffffff98000000680000006800000;
		6'b110101:	xpb = 256'h06a000000000000000000000069ffffffffffffff960000006a0000006a00000;
		6'b110110:	xpb = 256'h06c00000000000000000000006bffffffffffffff940000006c0000006c00000;
		6'b110111:	xpb = 256'h06e00000000000000000000006dffffffffffffff920000006e0000006e00000;
		6'b111000:	xpb = 256'h07000000000000000000000006fffffffffffffff90000000700000007000000;
		6'b111001:	xpb = 256'h072000000000000000000000071ffffffffffffff8e000000720000007200000;
		6'b111010:	xpb = 256'h074000000000000000000000073ffffffffffffff8c000000740000007400000;
		6'b111011:	xpb = 256'h076000000000000000000000075ffffffffffffff8a000000760000007600000;
		6'b111100:	xpb = 256'h078000000000000000000000077ffffffffffffff88000000780000007800000;
		6'b111101:	xpb = 256'h07a000000000000000000000079ffffffffffffff860000007a0000007a00000;
		6'b111110:	xpb = 256'h07c00000000000000000000007bffffffffffffff840000007c0000007c00000;
		6'b111111:	xpb = 256'h07e00000000000000000000007dffffffffffffff820000007e0000007e00000;
	endcase
end
endmodule

module xpb_19_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h08000000000000000000000007fffffffffffffff80000000800000008000000;
		6'b000010:	xpb = 256'h1000000000000000000000000ffffffffffffffff00000001000000010000000;
		6'b000011:	xpb = 256'h18000000000000000000000017ffffffffffffffe80000001800000018000000;
		6'b000100:	xpb = 256'h2000000000000000000000001fffffffffffffffe00000002000000020000000;
		6'b000101:	xpb = 256'h28000000000000000000000027ffffffffffffffd80000002800000028000000;
		6'b000110:	xpb = 256'h3000000000000000000000002fffffffffffffffd00000003000000030000000;
		6'b000111:	xpb = 256'h38000000000000000000000037ffffffffffffffc80000003800000038000000;
		6'b001000:	xpb = 256'h4000000000000000000000003fffffffffffffffc00000004000000040000000;
		6'b001001:	xpb = 256'h48000000000000000000000047ffffffffffffffb80000004800000048000000;
		6'b001010:	xpb = 256'h5000000000000000000000004fffffffffffffffb00000005000000050000000;
		6'b001011:	xpb = 256'h58000000000000000000000057ffffffffffffffa80000005800000058000000;
		6'b001100:	xpb = 256'h6000000000000000000000005fffffffffffffffa00000006000000060000000;
		6'b001101:	xpb = 256'h68000000000000000000000067ffffffffffffff980000006800000068000000;
		6'b001110:	xpb = 256'h7000000000000000000000006fffffffffffffff900000007000000070000000;
		6'b001111:	xpb = 256'h78000000000000000000000077ffffffffffffff880000007800000078000000;
		6'b010000:	xpb = 256'h8000000000000000000000007fffffffffffffff800000008000000080000000;
		6'b010001:	xpb = 256'h88000000000000000000000087ffffffffffffff780000008800000088000000;
		6'b010010:	xpb = 256'h9000000000000000000000008fffffffffffffff700000009000000090000000;
		6'b010011:	xpb = 256'h98000000000000000000000097ffffffffffffff680000009800000098000000;
		6'b010100:	xpb = 256'ha000000000000000000000009fffffffffffffff60000000a0000000a0000000;
		6'b010101:	xpb = 256'ha80000000000000000000000a7ffffffffffffff58000000a8000000a8000000;
		6'b010110:	xpb = 256'hb00000000000000000000000afffffffffffffff50000000b0000000b0000000;
		6'b010111:	xpb = 256'hb80000000000000000000000b7ffffffffffffff48000000b8000000b8000000;
		6'b011000:	xpb = 256'hc00000000000000000000000bfffffffffffffff40000000c0000000c0000000;
		6'b011001:	xpb = 256'hc80000000000000000000000c7ffffffffffffff38000000c8000000c8000000;
		6'b011010:	xpb = 256'hd00000000000000000000000cfffffffffffffff30000000d0000000d0000000;
		6'b011011:	xpb = 256'hd80000000000000000000000d7ffffffffffffff28000000d8000000d8000000;
		6'b011100:	xpb = 256'he00000000000000000000000dfffffffffffffff20000000e0000000e0000000;
		6'b011101:	xpb = 256'he80000000000000000000000e7ffffffffffffff18000000e8000000e8000000;
		6'b011110:	xpb = 256'hf00000000000000000000000efffffffffffffff10000000f0000000f0000000;
		6'b011111:	xpb = 256'hf80000000000000000000000f7ffffffffffffff08000000f8000000f8000000;
		6'b100000:	xpb = 256'h0000000100000000000000010000000000000000000000000000000100000001;
		6'b100001:	xpb = 256'h08000001000000000000000107fffffffffffffff80000000800000108000001;
		6'b100010:	xpb = 256'h1000000100000000000000010ffffffffffffffff00000001000000110000001;
		6'b100011:	xpb = 256'h18000001000000000000000117ffffffffffffffe80000001800000118000001;
		6'b100100:	xpb = 256'h2000000100000000000000011fffffffffffffffe00000002000000120000001;
		6'b100101:	xpb = 256'h28000001000000000000000127ffffffffffffffd80000002800000128000001;
		6'b100110:	xpb = 256'h3000000100000000000000012fffffffffffffffd00000003000000130000001;
		6'b100111:	xpb = 256'h38000001000000000000000137ffffffffffffffc80000003800000138000001;
		6'b101000:	xpb = 256'h4000000100000000000000013fffffffffffffffc00000004000000140000001;
		6'b101001:	xpb = 256'h48000001000000000000000147ffffffffffffffb80000004800000148000001;
		6'b101010:	xpb = 256'h5000000100000000000000014fffffffffffffffb00000005000000150000001;
		6'b101011:	xpb = 256'h58000001000000000000000157ffffffffffffffa80000005800000158000001;
		6'b101100:	xpb = 256'h6000000100000000000000015fffffffffffffffa00000006000000160000001;
		6'b101101:	xpb = 256'h68000001000000000000000167ffffffffffffff980000006800000168000001;
		6'b101110:	xpb = 256'h7000000100000000000000016fffffffffffffff900000007000000170000001;
		6'b101111:	xpb = 256'h78000001000000000000000177ffffffffffffff880000007800000178000001;
		6'b110000:	xpb = 256'h8000000100000000000000017fffffffffffffff800000008000000180000001;
		6'b110001:	xpb = 256'h88000001000000000000000187ffffffffffffff780000008800000188000001;
		6'b110010:	xpb = 256'h9000000100000000000000018fffffffffffffff700000009000000190000001;
		6'b110011:	xpb = 256'h98000001000000000000000197ffffffffffffff680000009800000198000001;
		6'b110100:	xpb = 256'ha000000100000000000000019fffffffffffffff60000000a0000001a0000001;
		6'b110101:	xpb = 256'ha80000010000000000000001a7ffffffffffffff58000000a8000001a8000001;
		6'b110110:	xpb = 256'hb00000010000000000000001afffffffffffffff50000000b0000001b0000001;
		6'b110111:	xpb = 256'hb80000010000000000000001b7ffffffffffffff48000000b8000001b8000001;
		6'b111000:	xpb = 256'hc00000010000000000000001bfffffffffffffff40000000c0000001c0000001;
		6'b111001:	xpb = 256'hc80000010000000000000001c7ffffffffffffff38000000c8000001c8000001;
		6'b111010:	xpb = 256'hd00000010000000000000001cfffffffffffffff30000000d0000001d0000001;
		6'b111011:	xpb = 256'hd80000010000000000000001d7ffffffffffffff28000000d8000001d8000001;
		6'b111100:	xpb = 256'he00000010000000000000001dfffffffffffffff20000000e0000001e0000001;
		6'b111101:	xpb = 256'he80000010000000000000001e7ffffffffffffff18000000e8000001e8000001;
		6'b111110:	xpb = 256'hf00000010000000000000001efffffffffffffff10000000f0000001f0000001;
		6'b111111:	xpb = 256'hf80000010000000000000001f7ffffffffffffff08000000f8000001f8000001;
	endcase
end
endmodule

module xpb_20_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000100000000000000010000000000000000000000000000000100000001;
		5'b00010:	xpb = 256'h0000000200000000000000020000000000000000000000000000000200000002;
		5'b00011:	xpb = 256'h0000000300000000000000030000000000000000000000000000000300000003;
		5'b00100:	xpb = 256'h0000000400000000000000040000000000000000000000000000000400000004;
		5'b00101:	xpb = 256'h0000000500000000000000050000000000000000000000000000000500000005;
		5'b00110:	xpb = 256'h0000000600000000000000060000000000000000000000000000000600000006;
		5'b00111:	xpb = 256'h0000000700000000000000070000000000000000000000000000000700000007;
		5'b01000:	xpb = 256'h0000000800000000000000080000000000000000000000000000000800000008;
		5'b01001:	xpb = 256'h0000000900000000000000090000000000000000000000000000000900000009;
		5'b01010:	xpb = 256'h0000000a000000000000000a0000000000000000000000000000000a0000000a;
		5'b01011:	xpb = 256'h0000000b000000000000000b0000000000000000000000000000000b0000000b;
		5'b01100:	xpb = 256'h0000000c000000000000000c0000000000000000000000000000000c0000000c;
		5'b01101:	xpb = 256'h0000000d000000000000000d0000000000000000000000000000000d0000000d;
		5'b01110:	xpb = 256'h0000000e000000000000000e0000000000000000000000000000000e0000000e;
		5'b01111:	xpb = 256'h0000000f000000000000000f0000000000000000000000000000000f0000000f;
		5'b10000:	xpb = 256'h0000001000000000000000100000000000000000000000000000001000000010;
		5'b10001:	xpb = 256'h0000001100000000000000110000000000000000000000000000001100000011;
		5'b10010:	xpb = 256'h0000001200000000000000120000000000000000000000000000001200000012;
		5'b10011:	xpb = 256'h0000001300000000000000130000000000000000000000000000001300000013;
		5'b10100:	xpb = 256'h0000001400000000000000140000000000000000000000000000001400000014;
		5'b10101:	xpb = 256'h0000001500000000000000150000000000000000000000000000001500000015;
		5'b10110:	xpb = 256'h0000001600000000000000160000000000000000000000000000001600000016;
		5'b10111:	xpb = 256'h0000001700000000000000170000000000000000000000000000001700000017;
		5'b11000:	xpb = 256'h0000001800000000000000180000000000000000000000000000001800000018;
		5'b11001:	xpb = 256'h0000001900000000000000190000000000000000000000000000001900000019;
		5'b11010:	xpb = 256'h0000001a000000000000001a0000000000000000000000000000001a0000001a;
		5'b11011:	xpb = 256'h0000001b000000000000001b0000000000000000000000000000001b0000001b;
		5'b11100:	xpb = 256'h0000001c000000000000001c0000000000000000000000000000001c0000001c;
		5'b11101:	xpb = 256'h0000001d000000000000001d0000000000000000000000000000001d0000001d;
		5'b11110:	xpb = 256'h0000001e000000000000001e0000000000000000000000000000001e0000001e;
		5'b11111:	xpb = 256'h0000001f000000000000001f0000000000000000000000000000001f0000001f;
	endcase
end
endmodule

module xpb_20_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000002000000000000000200000000000000000000000000000002000000020;
		6'b000010:	xpb = 256'h0000004000000000000000400000000000000000000000000000004000000040;
		6'b000011:	xpb = 256'h0000006000000000000000600000000000000000000000000000006000000060;
		6'b000100:	xpb = 256'h0000008000000000000000800000000000000000000000000000008000000080;
		6'b000101:	xpb = 256'h000000a000000000000000a0000000000000000000000000000000a0000000a0;
		6'b000110:	xpb = 256'h000000c000000000000000c0000000000000000000000000000000c0000000c0;
		6'b000111:	xpb = 256'h000000e000000000000000e0000000000000000000000000000000e0000000e0;
		6'b001000:	xpb = 256'h0000010000000000000001000000000000000000000000000000010000000100;
		6'b001001:	xpb = 256'h0000012000000000000001200000000000000000000000000000012000000120;
		6'b001010:	xpb = 256'h0000014000000000000001400000000000000000000000000000014000000140;
		6'b001011:	xpb = 256'h0000016000000000000001600000000000000000000000000000016000000160;
		6'b001100:	xpb = 256'h0000018000000000000001800000000000000000000000000000018000000180;
		6'b001101:	xpb = 256'h000001a000000000000001a0000000000000000000000000000001a0000001a0;
		6'b001110:	xpb = 256'h000001c000000000000001c0000000000000000000000000000001c0000001c0;
		6'b001111:	xpb = 256'h000001e000000000000001e0000000000000000000000000000001e0000001e0;
		6'b010000:	xpb = 256'h0000020000000000000002000000000000000000000000000000020000000200;
		6'b010001:	xpb = 256'h0000022000000000000002200000000000000000000000000000022000000220;
		6'b010010:	xpb = 256'h0000024000000000000002400000000000000000000000000000024000000240;
		6'b010011:	xpb = 256'h0000026000000000000002600000000000000000000000000000026000000260;
		6'b010100:	xpb = 256'h0000028000000000000002800000000000000000000000000000028000000280;
		6'b010101:	xpb = 256'h000002a000000000000002a0000000000000000000000000000002a0000002a0;
		6'b010110:	xpb = 256'h000002c000000000000002c0000000000000000000000000000002c0000002c0;
		6'b010111:	xpb = 256'h000002e000000000000002e0000000000000000000000000000002e0000002e0;
		6'b011000:	xpb = 256'h0000030000000000000003000000000000000000000000000000030000000300;
		6'b011001:	xpb = 256'h0000032000000000000003200000000000000000000000000000032000000320;
		6'b011010:	xpb = 256'h0000034000000000000003400000000000000000000000000000034000000340;
		6'b011011:	xpb = 256'h0000036000000000000003600000000000000000000000000000036000000360;
		6'b011100:	xpb = 256'h0000038000000000000003800000000000000000000000000000038000000380;
		6'b011101:	xpb = 256'h000003a000000000000003a0000000000000000000000000000003a0000003a0;
		6'b011110:	xpb = 256'h000003c000000000000003c0000000000000000000000000000003c0000003c0;
		6'b011111:	xpb = 256'h000003e000000000000003e0000000000000000000000000000003e0000003e0;
		6'b100000:	xpb = 256'h0000040000000000000004000000000000000000000000000000040000000400;
		6'b100001:	xpb = 256'h0000042000000000000004200000000000000000000000000000042000000420;
		6'b100010:	xpb = 256'h0000044000000000000004400000000000000000000000000000044000000440;
		6'b100011:	xpb = 256'h0000046000000000000004600000000000000000000000000000046000000460;
		6'b100100:	xpb = 256'h0000048000000000000004800000000000000000000000000000048000000480;
		6'b100101:	xpb = 256'h000004a000000000000004a0000000000000000000000000000004a0000004a0;
		6'b100110:	xpb = 256'h000004c000000000000004c0000000000000000000000000000004c0000004c0;
		6'b100111:	xpb = 256'h000004e000000000000004e0000000000000000000000000000004e0000004e0;
		6'b101000:	xpb = 256'h0000050000000000000005000000000000000000000000000000050000000500;
		6'b101001:	xpb = 256'h0000052000000000000005200000000000000000000000000000052000000520;
		6'b101010:	xpb = 256'h0000054000000000000005400000000000000000000000000000054000000540;
		6'b101011:	xpb = 256'h0000056000000000000005600000000000000000000000000000056000000560;
		6'b101100:	xpb = 256'h0000058000000000000005800000000000000000000000000000058000000580;
		6'b101101:	xpb = 256'h000005a000000000000005a0000000000000000000000000000005a0000005a0;
		6'b101110:	xpb = 256'h000005c000000000000005c0000000000000000000000000000005c0000005c0;
		6'b101111:	xpb = 256'h000005e000000000000005e0000000000000000000000000000005e0000005e0;
		6'b110000:	xpb = 256'h0000060000000000000006000000000000000000000000000000060000000600;
		6'b110001:	xpb = 256'h0000062000000000000006200000000000000000000000000000062000000620;
		6'b110010:	xpb = 256'h0000064000000000000006400000000000000000000000000000064000000640;
		6'b110011:	xpb = 256'h0000066000000000000006600000000000000000000000000000066000000660;
		6'b110100:	xpb = 256'h0000068000000000000006800000000000000000000000000000068000000680;
		6'b110101:	xpb = 256'h000006a000000000000006a0000000000000000000000000000006a0000006a0;
		6'b110110:	xpb = 256'h000006c000000000000006c0000000000000000000000000000006c0000006c0;
		6'b110111:	xpb = 256'h000006e000000000000006e0000000000000000000000000000006e0000006e0;
		6'b111000:	xpb = 256'h0000070000000000000007000000000000000000000000000000070000000700;
		6'b111001:	xpb = 256'h0000072000000000000007200000000000000000000000000000072000000720;
		6'b111010:	xpb = 256'h0000074000000000000007400000000000000000000000000000074000000740;
		6'b111011:	xpb = 256'h0000076000000000000007600000000000000000000000000000076000000760;
		6'b111100:	xpb = 256'h0000078000000000000007800000000000000000000000000000078000000780;
		6'b111101:	xpb = 256'h000007a000000000000007a0000000000000000000000000000007a0000007a0;
		6'b111110:	xpb = 256'h000007c000000000000007c0000000000000000000000000000007c0000007c0;
		6'b111111:	xpb = 256'h000007e000000000000007e0000000000000000000000000000007e0000007e0;
	endcase
end
endmodule

module xpb_20_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000080000000000000008000000000000000000000000000000080000000800;
		6'b000010:	xpb = 256'h0000100000000000000010000000000000000000000000000000100000001000;
		6'b000011:	xpb = 256'h0000180000000000000018000000000000000000000000000000180000001800;
		6'b000100:	xpb = 256'h0000200000000000000020000000000000000000000000000000200000002000;
		6'b000101:	xpb = 256'h0000280000000000000028000000000000000000000000000000280000002800;
		6'b000110:	xpb = 256'h0000300000000000000030000000000000000000000000000000300000003000;
		6'b000111:	xpb = 256'h0000380000000000000038000000000000000000000000000000380000003800;
		6'b001000:	xpb = 256'h0000400000000000000040000000000000000000000000000000400000004000;
		6'b001001:	xpb = 256'h0000480000000000000048000000000000000000000000000000480000004800;
		6'b001010:	xpb = 256'h0000500000000000000050000000000000000000000000000000500000005000;
		6'b001011:	xpb = 256'h0000580000000000000058000000000000000000000000000000580000005800;
		6'b001100:	xpb = 256'h0000600000000000000060000000000000000000000000000000600000006000;
		6'b001101:	xpb = 256'h0000680000000000000068000000000000000000000000000000680000006800;
		6'b001110:	xpb = 256'h0000700000000000000070000000000000000000000000000000700000007000;
		6'b001111:	xpb = 256'h0000780000000000000078000000000000000000000000000000780000007800;
		6'b010000:	xpb = 256'h0000800000000000000080000000000000000000000000000000800000008000;
		6'b010001:	xpb = 256'h0000880000000000000088000000000000000000000000000000880000008800;
		6'b010010:	xpb = 256'h0000900000000000000090000000000000000000000000000000900000009000;
		6'b010011:	xpb = 256'h0000980000000000000098000000000000000000000000000000980000009800;
		6'b010100:	xpb = 256'h0000a000000000000000a0000000000000000000000000000000a0000000a000;
		6'b010101:	xpb = 256'h0000a800000000000000a8000000000000000000000000000000a8000000a800;
		6'b010110:	xpb = 256'h0000b000000000000000b0000000000000000000000000000000b0000000b000;
		6'b010111:	xpb = 256'h0000b800000000000000b8000000000000000000000000000000b8000000b800;
		6'b011000:	xpb = 256'h0000c000000000000000c0000000000000000000000000000000c0000000c000;
		6'b011001:	xpb = 256'h0000c800000000000000c8000000000000000000000000000000c8000000c800;
		6'b011010:	xpb = 256'h0000d000000000000000d0000000000000000000000000000000d0000000d000;
		6'b011011:	xpb = 256'h0000d800000000000000d8000000000000000000000000000000d8000000d800;
		6'b011100:	xpb = 256'h0000e000000000000000e0000000000000000000000000000000e0000000e000;
		6'b011101:	xpb = 256'h0000e800000000000000e8000000000000000000000000000000e8000000e800;
		6'b011110:	xpb = 256'h0000f000000000000000f0000000000000000000000000000000f0000000f000;
		6'b011111:	xpb = 256'h0000f800000000000000f8000000000000000000000000000000f8000000f800;
		6'b100000:	xpb = 256'h0001000000000000000100000000000000000000000000000001000000010000;
		6'b100001:	xpb = 256'h0001080000000000000108000000000000000000000000000001080000010800;
		6'b100010:	xpb = 256'h0001100000000000000110000000000000000000000000000001100000011000;
		6'b100011:	xpb = 256'h0001180000000000000118000000000000000000000000000001180000011800;
		6'b100100:	xpb = 256'h0001200000000000000120000000000000000000000000000001200000012000;
		6'b100101:	xpb = 256'h0001280000000000000128000000000000000000000000000001280000012800;
		6'b100110:	xpb = 256'h0001300000000000000130000000000000000000000000000001300000013000;
		6'b100111:	xpb = 256'h0001380000000000000138000000000000000000000000000001380000013800;
		6'b101000:	xpb = 256'h0001400000000000000140000000000000000000000000000001400000014000;
		6'b101001:	xpb = 256'h0001480000000000000148000000000000000000000000000001480000014800;
		6'b101010:	xpb = 256'h0001500000000000000150000000000000000000000000000001500000015000;
		6'b101011:	xpb = 256'h0001580000000000000158000000000000000000000000000001580000015800;
		6'b101100:	xpb = 256'h0001600000000000000160000000000000000000000000000001600000016000;
		6'b101101:	xpb = 256'h0001680000000000000168000000000000000000000000000001680000016800;
		6'b101110:	xpb = 256'h0001700000000000000170000000000000000000000000000001700000017000;
		6'b101111:	xpb = 256'h0001780000000000000178000000000000000000000000000001780000017800;
		6'b110000:	xpb = 256'h0001800000000000000180000000000000000000000000000001800000018000;
		6'b110001:	xpb = 256'h0001880000000000000188000000000000000000000000000001880000018800;
		6'b110010:	xpb = 256'h0001900000000000000190000000000000000000000000000001900000019000;
		6'b110011:	xpb = 256'h0001980000000000000198000000000000000000000000000001980000019800;
		6'b110100:	xpb = 256'h0001a000000000000001a0000000000000000000000000000001a0000001a000;
		6'b110101:	xpb = 256'h0001a800000000000001a8000000000000000000000000000001a8000001a800;
		6'b110110:	xpb = 256'h0001b000000000000001b0000000000000000000000000000001b0000001b000;
		6'b110111:	xpb = 256'h0001b800000000000001b8000000000000000000000000000001b8000001b800;
		6'b111000:	xpb = 256'h0001c000000000000001c0000000000000000000000000000001c0000001c000;
		6'b111001:	xpb = 256'h0001c800000000000001c8000000000000000000000000000001c8000001c800;
		6'b111010:	xpb = 256'h0001d000000000000001d0000000000000000000000000000001d0000001d000;
		6'b111011:	xpb = 256'h0001d800000000000001d8000000000000000000000000000001d8000001d800;
		6'b111100:	xpb = 256'h0001e000000000000001e0000000000000000000000000000001e0000001e000;
		6'b111101:	xpb = 256'h0001e800000000000001e8000000000000000000000000000001e8000001e800;
		6'b111110:	xpb = 256'h0001f000000000000001f0000000000000000000000000000001f0000001f000;
		6'b111111:	xpb = 256'h0001f800000000000001f8000000000000000000000000000001f8000001f800;
	endcase
end
endmodule

module xpb_21_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0001000000000000000100000000000000000000000000000001000000010000;
		5'b00010:	xpb = 256'h0002000000000000000200000000000000000000000000000002000000020000;
		5'b00011:	xpb = 256'h0003000000000000000300000000000000000000000000000003000000030000;
		5'b00100:	xpb = 256'h0004000000000000000400000000000000000000000000000004000000040000;
		5'b00101:	xpb = 256'h0005000000000000000500000000000000000000000000000005000000050000;
		5'b00110:	xpb = 256'h0006000000000000000600000000000000000000000000000006000000060000;
		5'b00111:	xpb = 256'h0007000000000000000700000000000000000000000000000007000000070000;
		5'b01000:	xpb = 256'h0008000000000000000800000000000000000000000000000008000000080000;
		5'b01001:	xpb = 256'h0009000000000000000900000000000000000000000000000009000000090000;
		5'b01010:	xpb = 256'h000a000000000000000a0000000000000000000000000000000a0000000a0000;
		5'b01011:	xpb = 256'h000b000000000000000b0000000000000000000000000000000b0000000b0000;
		5'b01100:	xpb = 256'h000c000000000000000c0000000000000000000000000000000c0000000c0000;
		5'b01101:	xpb = 256'h000d000000000000000d0000000000000000000000000000000d0000000d0000;
		5'b01110:	xpb = 256'h000e000000000000000e0000000000000000000000000000000e0000000e0000;
		5'b01111:	xpb = 256'h000f000000000000000f0000000000000000000000000000000f0000000f0000;
		5'b10000:	xpb = 256'h0010000000000000001000000000000000000000000000000010000000100000;
		5'b10001:	xpb = 256'h0011000000000000001100000000000000000000000000000011000000110000;
		5'b10010:	xpb = 256'h0012000000000000001200000000000000000000000000000012000000120000;
		5'b10011:	xpb = 256'h0013000000000000001300000000000000000000000000000013000000130000;
		5'b10100:	xpb = 256'h0014000000000000001400000000000000000000000000000014000000140000;
		5'b10101:	xpb = 256'h0015000000000000001500000000000000000000000000000015000000150000;
		5'b10110:	xpb = 256'h0016000000000000001600000000000000000000000000000016000000160000;
		5'b10111:	xpb = 256'h0017000000000000001700000000000000000000000000000017000000170000;
		5'b11000:	xpb = 256'h0018000000000000001800000000000000000000000000000018000000180000;
		5'b11001:	xpb = 256'h0019000000000000001900000000000000000000000000000019000000190000;
		5'b11010:	xpb = 256'h001a000000000000001a0000000000000000000000000000001a0000001a0000;
		5'b11011:	xpb = 256'h001b000000000000001b0000000000000000000000000000001b0000001b0000;
		5'b11100:	xpb = 256'h001c000000000000001c0000000000000000000000000000001c0000001c0000;
		5'b11101:	xpb = 256'h001d000000000000001d0000000000000000000000000000001d0000001d0000;
		5'b11110:	xpb = 256'h001e000000000000001e0000000000000000000000000000001e0000001e0000;
		5'b11111:	xpb = 256'h001f000000000000001f0000000000000000000000000000001f0000001f0000;
	endcase
end
endmodule

module xpb_21_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0020000000000000002000000000000000000000000000000020000000200000;
		6'b000010:	xpb = 256'h0040000000000000004000000000000000000000000000000040000000400000;
		6'b000011:	xpb = 256'h0060000000000000006000000000000000000000000000000060000000600000;
		6'b000100:	xpb = 256'h0080000000000000008000000000000000000000000000000080000000800000;
		6'b000101:	xpb = 256'h00a000000000000000a0000000000000000000000000000000a0000000a00000;
		6'b000110:	xpb = 256'h00c000000000000000c0000000000000000000000000000000c0000000c00000;
		6'b000111:	xpb = 256'h00e000000000000000e0000000000000000000000000000000e0000000e00000;
		6'b001000:	xpb = 256'h0100000000000000010000000000000000000000000000000100000001000000;
		6'b001001:	xpb = 256'h0120000000000000012000000000000000000000000000000120000001200000;
		6'b001010:	xpb = 256'h0140000000000000014000000000000000000000000000000140000001400000;
		6'b001011:	xpb = 256'h0160000000000000016000000000000000000000000000000160000001600000;
		6'b001100:	xpb = 256'h0180000000000000018000000000000000000000000000000180000001800000;
		6'b001101:	xpb = 256'h01a000000000000001a0000000000000000000000000000001a0000001a00000;
		6'b001110:	xpb = 256'h01c000000000000001c0000000000000000000000000000001c0000001c00000;
		6'b001111:	xpb = 256'h01e000000000000001e0000000000000000000000000000001e0000001e00000;
		6'b010000:	xpb = 256'h0200000000000000020000000000000000000000000000000200000002000000;
		6'b010001:	xpb = 256'h0220000000000000022000000000000000000000000000000220000002200000;
		6'b010010:	xpb = 256'h0240000000000000024000000000000000000000000000000240000002400000;
		6'b010011:	xpb = 256'h0260000000000000026000000000000000000000000000000260000002600000;
		6'b010100:	xpb = 256'h0280000000000000028000000000000000000000000000000280000002800000;
		6'b010101:	xpb = 256'h02a000000000000002a0000000000000000000000000000002a0000002a00000;
		6'b010110:	xpb = 256'h02c000000000000002c0000000000000000000000000000002c0000002c00000;
		6'b010111:	xpb = 256'h02e000000000000002e0000000000000000000000000000002e0000002e00000;
		6'b011000:	xpb = 256'h0300000000000000030000000000000000000000000000000300000003000000;
		6'b011001:	xpb = 256'h0320000000000000032000000000000000000000000000000320000003200000;
		6'b011010:	xpb = 256'h0340000000000000034000000000000000000000000000000340000003400000;
		6'b011011:	xpb = 256'h0360000000000000036000000000000000000000000000000360000003600000;
		6'b011100:	xpb = 256'h0380000000000000038000000000000000000000000000000380000003800000;
		6'b011101:	xpb = 256'h03a000000000000003a0000000000000000000000000000003a0000003a00000;
		6'b011110:	xpb = 256'h03c000000000000003c0000000000000000000000000000003c0000003c00000;
		6'b011111:	xpb = 256'h03e000000000000003e0000000000000000000000000000003e0000003e00000;
		6'b100000:	xpb = 256'h0400000000000000040000000000000000000000000000000400000004000000;
		6'b100001:	xpb = 256'h0420000000000000042000000000000000000000000000000420000004200000;
		6'b100010:	xpb = 256'h0440000000000000044000000000000000000000000000000440000004400000;
		6'b100011:	xpb = 256'h0460000000000000046000000000000000000000000000000460000004600000;
		6'b100100:	xpb = 256'h0480000000000000048000000000000000000000000000000480000004800000;
		6'b100101:	xpb = 256'h04a000000000000004a0000000000000000000000000000004a0000004a00000;
		6'b100110:	xpb = 256'h04c000000000000004c0000000000000000000000000000004c0000004c00000;
		6'b100111:	xpb = 256'h04e000000000000004e0000000000000000000000000000004e0000004e00000;
		6'b101000:	xpb = 256'h0500000000000000050000000000000000000000000000000500000005000000;
		6'b101001:	xpb = 256'h0520000000000000052000000000000000000000000000000520000005200000;
		6'b101010:	xpb = 256'h0540000000000000054000000000000000000000000000000540000005400000;
		6'b101011:	xpb = 256'h0560000000000000056000000000000000000000000000000560000005600000;
		6'b101100:	xpb = 256'h0580000000000000058000000000000000000000000000000580000005800000;
		6'b101101:	xpb = 256'h05a000000000000005a0000000000000000000000000000005a0000005a00000;
		6'b101110:	xpb = 256'h05c000000000000005c0000000000000000000000000000005c0000005c00000;
		6'b101111:	xpb = 256'h05e000000000000005e0000000000000000000000000000005e0000005e00000;
		6'b110000:	xpb = 256'h0600000000000000060000000000000000000000000000000600000006000000;
		6'b110001:	xpb = 256'h0620000000000000062000000000000000000000000000000620000006200000;
		6'b110010:	xpb = 256'h0640000000000000064000000000000000000000000000000640000006400000;
		6'b110011:	xpb = 256'h0660000000000000066000000000000000000000000000000660000006600000;
		6'b110100:	xpb = 256'h0680000000000000068000000000000000000000000000000680000006800000;
		6'b110101:	xpb = 256'h06a000000000000006a0000000000000000000000000000006a0000006a00000;
		6'b110110:	xpb = 256'h06c000000000000006c0000000000000000000000000000006c0000006c00000;
		6'b110111:	xpb = 256'h06e000000000000006e0000000000000000000000000000006e0000006e00000;
		6'b111000:	xpb = 256'h0700000000000000070000000000000000000000000000000700000007000000;
		6'b111001:	xpb = 256'h0720000000000000072000000000000000000000000000000720000007200000;
		6'b111010:	xpb = 256'h0740000000000000074000000000000000000000000000000740000007400000;
		6'b111011:	xpb = 256'h0760000000000000076000000000000000000000000000000760000007600000;
		6'b111100:	xpb = 256'h0780000000000000078000000000000000000000000000000780000007800000;
		6'b111101:	xpb = 256'h07a000000000000007a0000000000000000000000000000007a0000007a00000;
		6'b111110:	xpb = 256'h07c000000000000007c0000000000000000000000000000007c0000007c00000;
		6'b111111:	xpb = 256'h07e000000000000007e0000000000000000000000000000007e0000007e00000;
	endcase
end
endmodule

module xpb_21_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0800000000000000080000000000000000000000000000000800000008000000;
		6'b000010:	xpb = 256'h1000000000000000100000000000000000000000000000001000000010000000;
		6'b000011:	xpb = 256'h1800000000000000180000000000000000000000000000001800000018000000;
		6'b000100:	xpb = 256'h2000000000000000200000000000000000000000000000002000000020000000;
		6'b000101:	xpb = 256'h2800000000000000280000000000000000000000000000002800000028000000;
		6'b000110:	xpb = 256'h3000000000000000300000000000000000000000000000003000000030000000;
		6'b000111:	xpb = 256'h3800000000000000380000000000000000000000000000003800000038000000;
		6'b001000:	xpb = 256'h4000000000000000400000000000000000000000000000004000000040000000;
		6'b001001:	xpb = 256'h4800000000000000480000000000000000000000000000004800000048000000;
		6'b001010:	xpb = 256'h5000000000000000500000000000000000000000000000005000000050000000;
		6'b001011:	xpb = 256'h5800000000000000580000000000000000000000000000005800000058000000;
		6'b001100:	xpb = 256'h6000000000000000600000000000000000000000000000006000000060000000;
		6'b001101:	xpb = 256'h6800000000000000680000000000000000000000000000006800000068000000;
		6'b001110:	xpb = 256'h7000000000000000700000000000000000000000000000007000000070000000;
		6'b001111:	xpb = 256'h7800000000000000780000000000000000000000000000007800000078000000;
		6'b010000:	xpb = 256'h8000000000000000800000000000000000000000000000008000000080000000;
		6'b010001:	xpb = 256'h8800000000000000880000000000000000000000000000008800000088000000;
		6'b010010:	xpb = 256'h9000000000000000900000000000000000000000000000009000000090000000;
		6'b010011:	xpb = 256'h9800000000000000980000000000000000000000000000009800000098000000;
		6'b010100:	xpb = 256'ha000000000000000a0000000000000000000000000000000a0000000a0000000;
		6'b010101:	xpb = 256'ha800000000000000a8000000000000000000000000000000a8000000a8000000;
		6'b010110:	xpb = 256'hb000000000000000b0000000000000000000000000000000b0000000b0000000;
		6'b010111:	xpb = 256'hb800000000000000b8000000000000000000000000000000b8000000b8000000;
		6'b011000:	xpb = 256'hc000000000000000c0000000000000000000000000000000c0000000c0000000;
		6'b011001:	xpb = 256'hc800000000000000c8000000000000000000000000000000c8000000c8000000;
		6'b011010:	xpb = 256'hd000000000000000d0000000000000000000000000000000d0000000d0000000;
		6'b011011:	xpb = 256'hd800000000000000d8000000000000000000000000000000d8000000d8000000;
		6'b011100:	xpb = 256'he000000000000000e0000000000000000000000000000000e0000000e0000000;
		6'b011101:	xpb = 256'he800000000000000e8000000000000000000000000000000e8000000e8000000;
		6'b011110:	xpb = 256'hf000000000000000f0000000000000000000000000000000f0000000f0000000;
		6'b011111:	xpb = 256'hf800000000000000f8000000000000000000000000000000f8000000f8000000;
		6'b100000:	xpb = 256'h0000000100000001000000000000000000000001000000000000000100000001;
		6'b100001:	xpb = 256'h0800000100000001080000000000000000000001000000000800000108000001;
		6'b100010:	xpb = 256'h1000000100000001100000000000000000000001000000001000000110000001;
		6'b100011:	xpb = 256'h1800000100000001180000000000000000000001000000001800000118000001;
		6'b100100:	xpb = 256'h2000000100000001200000000000000000000001000000002000000120000001;
		6'b100101:	xpb = 256'h2800000100000001280000000000000000000001000000002800000128000001;
		6'b100110:	xpb = 256'h3000000100000001300000000000000000000001000000003000000130000001;
		6'b100111:	xpb = 256'h3800000100000001380000000000000000000001000000003800000138000001;
		6'b101000:	xpb = 256'h4000000100000001400000000000000000000001000000004000000140000001;
		6'b101001:	xpb = 256'h4800000100000001480000000000000000000001000000004800000148000001;
		6'b101010:	xpb = 256'h5000000100000001500000000000000000000001000000005000000150000001;
		6'b101011:	xpb = 256'h5800000100000001580000000000000000000001000000005800000158000001;
		6'b101100:	xpb = 256'h6000000100000001600000000000000000000001000000006000000160000001;
		6'b101101:	xpb = 256'h6800000100000001680000000000000000000001000000006800000168000001;
		6'b101110:	xpb = 256'h7000000100000001700000000000000000000001000000007000000170000001;
		6'b101111:	xpb = 256'h7800000100000001780000000000000000000001000000007800000178000001;
		6'b110000:	xpb = 256'h8000000100000001800000000000000000000001000000008000000180000001;
		6'b110001:	xpb = 256'h8800000100000001880000000000000000000001000000008800000188000001;
		6'b110010:	xpb = 256'h9000000100000001900000000000000000000001000000009000000190000001;
		6'b110011:	xpb = 256'h9800000100000001980000000000000000000001000000009800000198000001;
		6'b110100:	xpb = 256'ha000000100000001a0000000000000000000000100000000a0000001a0000001;
		6'b110101:	xpb = 256'ha800000100000001a8000000000000000000000100000000a8000001a8000001;
		6'b110110:	xpb = 256'hb000000100000001b0000000000000000000000100000000b0000001b0000001;
		6'b110111:	xpb = 256'hb800000100000001b8000000000000000000000100000000b8000001b8000001;
		6'b111000:	xpb = 256'hc000000100000001c0000000000000000000000100000000c0000001c0000001;
		6'b111001:	xpb = 256'hc800000100000001c8000000000000000000000100000000c8000001c8000001;
		6'b111010:	xpb = 256'hd000000100000001d0000000000000000000000100000000d0000001d0000001;
		6'b111011:	xpb = 256'hd800000100000001d8000000000000000000000100000000d8000001d8000001;
		6'b111100:	xpb = 256'he000000100000001e0000000000000000000000100000000e0000001e0000001;
		6'b111101:	xpb = 256'he800000100000001e8000000000000000000000100000000e8000001e8000001;
		6'b111110:	xpb = 256'hf000000100000001f0000000000000000000000100000000f0000001f0000001;
		6'b111111:	xpb = 256'hf800000100000001f8000000000000000000000100000000f8000001f8000001;
	endcase
end
endmodule

module xpb_22_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000100000001000000000000000000000001000000000000000100000001;
		5'b00010:	xpb = 256'h0000000200000002000000000000000000000002000000000000000200000002;
		5'b00011:	xpb = 256'h0000000300000003000000000000000000000003000000000000000300000003;
		5'b00100:	xpb = 256'h0000000400000004000000000000000000000004000000000000000400000004;
		5'b00101:	xpb = 256'h0000000500000005000000000000000000000005000000000000000500000005;
		5'b00110:	xpb = 256'h0000000600000006000000000000000000000006000000000000000600000006;
		5'b00111:	xpb = 256'h0000000700000007000000000000000000000007000000000000000700000007;
		5'b01000:	xpb = 256'h0000000800000008000000000000000000000008000000000000000800000008;
		5'b01001:	xpb = 256'h0000000900000009000000000000000000000009000000000000000900000009;
		5'b01010:	xpb = 256'h0000000a0000000a00000000000000000000000a000000000000000a0000000a;
		5'b01011:	xpb = 256'h0000000b0000000b00000000000000000000000b000000000000000b0000000b;
		5'b01100:	xpb = 256'h0000000c0000000c00000000000000000000000c000000000000000c0000000c;
		5'b01101:	xpb = 256'h0000000d0000000d00000000000000000000000d000000000000000d0000000d;
		5'b01110:	xpb = 256'h0000000e0000000e00000000000000000000000e000000000000000e0000000e;
		5'b01111:	xpb = 256'h0000000f0000000f00000000000000000000000f000000000000000f0000000f;
		5'b10000:	xpb = 256'h0000001000000010000000000000000000000010000000000000001000000010;
		5'b10001:	xpb = 256'h0000001100000011000000000000000000000011000000000000001100000011;
		5'b10010:	xpb = 256'h0000001200000012000000000000000000000012000000000000001200000012;
		5'b10011:	xpb = 256'h0000001300000013000000000000000000000013000000000000001300000013;
		5'b10100:	xpb = 256'h0000001400000014000000000000000000000014000000000000001400000014;
		5'b10101:	xpb = 256'h0000001500000015000000000000000000000015000000000000001500000015;
		5'b10110:	xpb = 256'h0000001600000016000000000000000000000016000000000000001600000016;
		5'b10111:	xpb = 256'h0000001700000017000000000000000000000017000000000000001700000017;
		5'b11000:	xpb = 256'h0000001800000018000000000000000000000018000000000000001800000018;
		5'b11001:	xpb = 256'h0000001900000019000000000000000000000019000000000000001900000019;
		5'b11010:	xpb = 256'h0000001a0000001a00000000000000000000001a000000000000001a0000001a;
		5'b11011:	xpb = 256'h0000001b0000001b00000000000000000000001b000000000000001b0000001b;
		5'b11100:	xpb = 256'h0000001c0000001c00000000000000000000001c000000000000001c0000001c;
		5'b11101:	xpb = 256'h0000001d0000001d00000000000000000000001d000000000000001d0000001d;
		5'b11110:	xpb = 256'h0000001e0000001e00000000000000000000001e000000000000001e0000001e;
		5'b11111:	xpb = 256'h0000001f0000001f00000000000000000000001f000000000000001f0000001f;
	endcase
end
endmodule

module xpb_22_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000002000000020000000000000000000000020000000000000002000000020;
		6'b000010:	xpb = 256'h0000004000000040000000000000000000000040000000000000004000000040;
		6'b000011:	xpb = 256'h0000006000000060000000000000000000000060000000000000006000000060;
		6'b000100:	xpb = 256'h0000008000000080000000000000000000000080000000000000008000000080;
		6'b000101:	xpb = 256'h000000a0000000a00000000000000000000000a000000000000000a0000000a0;
		6'b000110:	xpb = 256'h000000c0000000c00000000000000000000000c000000000000000c0000000c0;
		6'b000111:	xpb = 256'h000000e0000000e00000000000000000000000e000000000000000e0000000e0;
		6'b001000:	xpb = 256'h0000010000000100000000000000000000000100000000000000010000000100;
		6'b001001:	xpb = 256'h0000012000000120000000000000000000000120000000000000012000000120;
		6'b001010:	xpb = 256'h0000014000000140000000000000000000000140000000000000014000000140;
		6'b001011:	xpb = 256'h0000016000000160000000000000000000000160000000000000016000000160;
		6'b001100:	xpb = 256'h0000018000000180000000000000000000000180000000000000018000000180;
		6'b001101:	xpb = 256'h000001a0000001a00000000000000000000001a000000000000001a0000001a0;
		6'b001110:	xpb = 256'h000001c0000001c00000000000000000000001c000000000000001c0000001c0;
		6'b001111:	xpb = 256'h000001e0000001e00000000000000000000001e000000000000001e0000001e0;
		6'b010000:	xpb = 256'h0000020000000200000000000000000000000200000000000000020000000200;
		6'b010001:	xpb = 256'h0000022000000220000000000000000000000220000000000000022000000220;
		6'b010010:	xpb = 256'h0000024000000240000000000000000000000240000000000000024000000240;
		6'b010011:	xpb = 256'h0000026000000260000000000000000000000260000000000000026000000260;
		6'b010100:	xpb = 256'h0000028000000280000000000000000000000280000000000000028000000280;
		6'b010101:	xpb = 256'h000002a0000002a00000000000000000000002a000000000000002a0000002a0;
		6'b010110:	xpb = 256'h000002c0000002c00000000000000000000002c000000000000002c0000002c0;
		6'b010111:	xpb = 256'h000002e0000002e00000000000000000000002e000000000000002e0000002e0;
		6'b011000:	xpb = 256'h0000030000000300000000000000000000000300000000000000030000000300;
		6'b011001:	xpb = 256'h0000032000000320000000000000000000000320000000000000032000000320;
		6'b011010:	xpb = 256'h0000034000000340000000000000000000000340000000000000034000000340;
		6'b011011:	xpb = 256'h0000036000000360000000000000000000000360000000000000036000000360;
		6'b011100:	xpb = 256'h0000038000000380000000000000000000000380000000000000038000000380;
		6'b011101:	xpb = 256'h000003a0000003a00000000000000000000003a000000000000003a0000003a0;
		6'b011110:	xpb = 256'h000003c0000003c00000000000000000000003c000000000000003c0000003c0;
		6'b011111:	xpb = 256'h000003e0000003e00000000000000000000003e000000000000003e0000003e0;
		6'b100000:	xpb = 256'h0000040000000400000000000000000000000400000000000000040000000400;
		6'b100001:	xpb = 256'h0000042000000420000000000000000000000420000000000000042000000420;
		6'b100010:	xpb = 256'h0000044000000440000000000000000000000440000000000000044000000440;
		6'b100011:	xpb = 256'h0000046000000460000000000000000000000460000000000000046000000460;
		6'b100100:	xpb = 256'h0000048000000480000000000000000000000480000000000000048000000480;
		6'b100101:	xpb = 256'h000004a0000004a00000000000000000000004a000000000000004a0000004a0;
		6'b100110:	xpb = 256'h000004c0000004c00000000000000000000004c000000000000004c0000004c0;
		6'b100111:	xpb = 256'h000004e0000004e00000000000000000000004e000000000000004e0000004e0;
		6'b101000:	xpb = 256'h0000050000000500000000000000000000000500000000000000050000000500;
		6'b101001:	xpb = 256'h0000052000000520000000000000000000000520000000000000052000000520;
		6'b101010:	xpb = 256'h0000054000000540000000000000000000000540000000000000054000000540;
		6'b101011:	xpb = 256'h0000056000000560000000000000000000000560000000000000056000000560;
		6'b101100:	xpb = 256'h0000058000000580000000000000000000000580000000000000058000000580;
		6'b101101:	xpb = 256'h000005a0000005a00000000000000000000005a000000000000005a0000005a0;
		6'b101110:	xpb = 256'h000005c0000005c00000000000000000000005c000000000000005c0000005c0;
		6'b101111:	xpb = 256'h000005e0000005e00000000000000000000005e000000000000005e0000005e0;
		6'b110000:	xpb = 256'h0000060000000600000000000000000000000600000000000000060000000600;
		6'b110001:	xpb = 256'h0000062000000620000000000000000000000620000000000000062000000620;
		6'b110010:	xpb = 256'h0000064000000640000000000000000000000640000000000000064000000640;
		6'b110011:	xpb = 256'h0000066000000660000000000000000000000660000000000000066000000660;
		6'b110100:	xpb = 256'h0000068000000680000000000000000000000680000000000000068000000680;
		6'b110101:	xpb = 256'h000006a0000006a00000000000000000000006a000000000000006a0000006a0;
		6'b110110:	xpb = 256'h000006c0000006c00000000000000000000006c000000000000006c0000006c0;
		6'b110111:	xpb = 256'h000006e0000006e00000000000000000000006e000000000000006e0000006e0;
		6'b111000:	xpb = 256'h0000070000000700000000000000000000000700000000000000070000000700;
		6'b111001:	xpb = 256'h0000072000000720000000000000000000000720000000000000072000000720;
		6'b111010:	xpb = 256'h0000074000000740000000000000000000000740000000000000074000000740;
		6'b111011:	xpb = 256'h0000076000000760000000000000000000000760000000000000076000000760;
		6'b111100:	xpb = 256'h0000078000000780000000000000000000000780000000000000078000000780;
		6'b111101:	xpb = 256'h000007a0000007a00000000000000000000007a000000000000007a0000007a0;
		6'b111110:	xpb = 256'h000007c0000007c00000000000000000000007c000000000000007c0000007c0;
		6'b111111:	xpb = 256'h000007e0000007e00000000000000000000007e000000000000007e0000007e0;
	endcase
end
endmodule

module xpb_22_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000080000000800000000000000000000000800000000000000080000000800;
		6'b000010:	xpb = 256'h0000100000001000000000000000000000001000000000000000100000001000;
		6'b000011:	xpb = 256'h0000180000001800000000000000000000001800000000000000180000001800;
		6'b000100:	xpb = 256'h0000200000002000000000000000000000002000000000000000200000002000;
		6'b000101:	xpb = 256'h0000280000002800000000000000000000002800000000000000280000002800;
		6'b000110:	xpb = 256'h0000300000003000000000000000000000003000000000000000300000003000;
		6'b000111:	xpb = 256'h0000380000003800000000000000000000003800000000000000380000003800;
		6'b001000:	xpb = 256'h0000400000004000000000000000000000004000000000000000400000004000;
		6'b001001:	xpb = 256'h0000480000004800000000000000000000004800000000000000480000004800;
		6'b001010:	xpb = 256'h0000500000005000000000000000000000005000000000000000500000005000;
		6'b001011:	xpb = 256'h0000580000005800000000000000000000005800000000000000580000005800;
		6'b001100:	xpb = 256'h0000600000006000000000000000000000006000000000000000600000006000;
		6'b001101:	xpb = 256'h0000680000006800000000000000000000006800000000000000680000006800;
		6'b001110:	xpb = 256'h0000700000007000000000000000000000007000000000000000700000007000;
		6'b001111:	xpb = 256'h0000780000007800000000000000000000007800000000000000780000007800;
		6'b010000:	xpb = 256'h0000800000008000000000000000000000008000000000000000800000008000;
		6'b010001:	xpb = 256'h0000880000008800000000000000000000008800000000000000880000008800;
		6'b010010:	xpb = 256'h0000900000009000000000000000000000009000000000000000900000009000;
		6'b010011:	xpb = 256'h0000980000009800000000000000000000009800000000000000980000009800;
		6'b010100:	xpb = 256'h0000a0000000a00000000000000000000000a000000000000000a0000000a000;
		6'b010101:	xpb = 256'h0000a8000000a80000000000000000000000a800000000000000a8000000a800;
		6'b010110:	xpb = 256'h0000b0000000b00000000000000000000000b000000000000000b0000000b000;
		6'b010111:	xpb = 256'h0000b8000000b80000000000000000000000b800000000000000b8000000b800;
		6'b011000:	xpb = 256'h0000c0000000c00000000000000000000000c000000000000000c0000000c000;
		6'b011001:	xpb = 256'h0000c8000000c80000000000000000000000c800000000000000c8000000c800;
		6'b011010:	xpb = 256'h0000d0000000d00000000000000000000000d000000000000000d0000000d000;
		6'b011011:	xpb = 256'h0000d8000000d80000000000000000000000d800000000000000d8000000d800;
		6'b011100:	xpb = 256'h0000e0000000e00000000000000000000000e000000000000000e0000000e000;
		6'b011101:	xpb = 256'h0000e8000000e80000000000000000000000e800000000000000e8000000e800;
		6'b011110:	xpb = 256'h0000f0000000f00000000000000000000000f000000000000000f0000000f000;
		6'b011111:	xpb = 256'h0000f8000000f80000000000000000000000f800000000000000f8000000f800;
		6'b100000:	xpb = 256'h0001000000010000000000000000000000010000000000000001000000010000;
		6'b100001:	xpb = 256'h0001080000010800000000000000000000010800000000000001080000010800;
		6'b100010:	xpb = 256'h0001100000011000000000000000000000011000000000000001100000011000;
		6'b100011:	xpb = 256'h0001180000011800000000000000000000011800000000000001180000011800;
		6'b100100:	xpb = 256'h0001200000012000000000000000000000012000000000000001200000012000;
		6'b100101:	xpb = 256'h0001280000012800000000000000000000012800000000000001280000012800;
		6'b100110:	xpb = 256'h0001300000013000000000000000000000013000000000000001300000013000;
		6'b100111:	xpb = 256'h0001380000013800000000000000000000013800000000000001380000013800;
		6'b101000:	xpb = 256'h0001400000014000000000000000000000014000000000000001400000014000;
		6'b101001:	xpb = 256'h0001480000014800000000000000000000014800000000000001480000014800;
		6'b101010:	xpb = 256'h0001500000015000000000000000000000015000000000000001500000015000;
		6'b101011:	xpb = 256'h0001580000015800000000000000000000015800000000000001580000015800;
		6'b101100:	xpb = 256'h0001600000016000000000000000000000016000000000000001600000016000;
		6'b101101:	xpb = 256'h0001680000016800000000000000000000016800000000000001680000016800;
		6'b101110:	xpb = 256'h0001700000017000000000000000000000017000000000000001700000017000;
		6'b101111:	xpb = 256'h0001780000017800000000000000000000017800000000000001780000017800;
		6'b110000:	xpb = 256'h0001800000018000000000000000000000018000000000000001800000018000;
		6'b110001:	xpb = 256'h0001880000018800000000000000000000018800000000000001880000018800;
		6'b110010:	xpb = 256'h0001900000019000000000000000000000019000000000000001900000019000;
		6'b110011:	xpb = 256'h0001980000019800000000000000000000019800000000000001980000019800;
		6'b110100:	xpb = 256'h0001a0000001a00000000000000000000001a000000000000001a0000001a000;
		6'b110101:	xpb = 256'h0001a8000001a80000000000000000000001a800000000000001a8000001a800;
		6'b110110:	xpb = 256'h0001b0000001b00000000000000000000001b000000000000001b0000001b000;
		6'b110111:	xpb = 256'h0001b8000001b80000000000000000000001b800000000000001b8000001b800;
		6'b111000:	xpb = 256'h0001c0000001c00000000000000000000001c000000000000001c0000001c000;
		6'b111001:	xpb = 256'h0001c8000001c80000000000000000000001c800000000000001c8000001c800;
		6'b111010:	xpb = 256'h0001d0000001d00000000000000000000001d000000000000001d0000001d000;
		6'b111011:	xpb = 256'h0001d8000001d80000000000000000000001d800000000000001d8000001d800;
		6'b111100:	xpb = 256'h0001e0000001e00000000000000000000001e000000000000001e0000001e000;
		6'b111101:	xpb = 256'h0001e8000001e80000000000000000000001e800000000000001e8000001e800;
		6'b111110:	xpb = 256'h0001f0000001f00000000000000000000001f000000000000001f0000001f000;
		6'b111111:	xpb = 256'h0001f8000001f80000000000000000000001f800000000000001f8000001f800;
	endcase
end
endmodule

module xpb_23_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0001000000010000000000000000000000010000000000000001000000010000;
		5'b00010:	xpb = 256'h0002000000020000000000000000000000020000000000000002000000020000;
		5'b00011:	xpb = 256'h0003000000030000000000000000000000030000000000000003000000030000;
		5'b00100:	xpb = 256'h0004000000040000000000000000000000040000000000000004000000040000;
		5'b00101:	xpb = 256'h0005000000050000000000000000000000050000000000000005000000050000;
		5'b00110:	xpb = 256'h0006000000060000000000000000000000060000000000000006000000060000;
		5'b00111:	xpb = 256'h0007000000070000000000000000000000070000000000000007000000070000;
		5'b01000:	xpb = 256'h0008000000080000000000000000000000080000000000000008000000080000;
		5'b01001:	xpb = 256'h0009000000090000000000000000000000090000000000000009000000090000;
		5'b01010:	xpb = 256'h000a0000000a00000000000000000000000a000000000000000a0000000a0000;
		5'b01011:	xpb = 256'h000b0000000b00000000000000000000000b000000000000000b0000000b0000;
		5'b01100:	xpb = 256'h000c0000000c00000000000000000000000c000000000000000c0000000c0000;
		5'b01101:	xpb = 256'h000d0000000d00000000000000000000000d000000000000000d0000000d0000;
		5'b01110:	xpb = 256'h000e0000000e00000000000000000000000e000000000000000e0000000e0000;
		5'b01111:	xpb = 256'h000f0000000f00000000000000000000000f000000000000000f0000000f0000;
		5'b10000:	xpb = 256'h0010000000100000000000000000000000100000000000000010000000100000;
		5'b10001:	xpb = 256'h0011000000110000000000000000000000110000000000000011000000110000;
		5'b10010:	xpb = 256'h0012000000120000000000000000000000120000000000000012000000120000;
		5'b10011:	xpb = 256'h0013000000130000000000000000000000130000000000000013000000130000;
		5'b10100:	xpb = 256'h0014000000140000000000000000000000140000000000000014000000140000;
		5'b10101:	xpb = 256'h0015000000150000000000000000000000150000000000000015000000150000;
		5'b10110:	xpb = 256'h0016000000160000000000000000000000160000000000000016000000160000;
		5'b10111:	xpb = 256'h0017000000170000000000000000000000170000000000000017000000170000;
		5'b11000:	xpb = 256'h0018000000180000000000000000000000180000000000000018000000180000;
		5'b11001:	xpb = 256'h0019000000190000000000000000000000190000000000000019000000190000;
		5'b11010:	xpb = 256'h001a0000001a00000000000000000000001a000000000000001a0000001a0000;
		5'b11011:	xpb = 256'h001b0000001b00000000000000000000001b000000000000001b0000001b0000;
		5'b11100:	xpb = 256'h001c0000001c00000000000000000000001c000000000000001c0000001c0000;
		5'b11101:	xpb = 256'h001d0000001d00000000000000000000001d000000000000001d0000001d0000;
		5'b11110:	xpb = 256'h001e0000001e00000000000000000000001e000000000000001e0000001e0000;
		5'b11111:	xpb = 256'h001f0000001f00000000000000000000001f000000000000001f0000001f0000;
	endcase
end
endmodule

module xpb_23_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0020000000200000000000000000000000200000000000000020000000200000;
		6'b000010:	xpb = 256'h0040000000400000000000000000000000400000000000000040000000400000;
		6'b000011:	xpb = 256'h0060000000600000000000000000000000600000000000000060000000600000;
		6'b000100:	xpb = 256'h0080000000800000000000000000000000800000000000000080000000800000;
		6'b000101:	xpb = 256'h00a0000000a00000000000000000000000a000000000000000a0000000a00000;
		6'b000110:	xpb = 256'h00c0000000c00000000000000000000000c000000000000000c0000000c00000;
		6'b000111:	xpb = 256'h00e0000000e00000000000000000000000e000000000000000e0000000e00000;
		6'b001000:	xpb = 256'h0100000001000000000000000000000001000000000000000100000001000000;
		6'b001001:	xpb = 256'h0120000001200000000000000000000001200000000000000120000001200000;
		6'b001010:	xpb = 256'h0140000001400000000000000000000001400000000000000140000001400000;
		6'b001011:	xpb = 256'h0160000001600000000000000000000001600000000000000160000001600000;
		6'b001100:	xpb = 256'h0180000001800000000000000000000001800000000000000180000001800000;
		6'b001101:	xpb = 256'h01a0000001a00000000000000000000001a000000000000001a0000001a00000;
		6'b001110:	xpb = 256'h01c0000001c00000000000000000000001c000000000000001c0000001c00000;
		6'b001111:	xpb = 256'h01e0000001e00000000000000000000001e000000000000001e0000001e00000;
		6'b010000:	xpb = 256'h0200000002000000000000000000000002000000000000000200000002000000;
		6'b010001:	xpb = 256'h0220000002200000000000000000000002200000000000000220000002200000;
		6'b010010:	xpb = 256'h0240000002400000000000000000000002400000000000000240000002400000;
		6'b010011:	xpb = 256'h0260000002600000000000000000000002600000000000000260000002600000;
		6'b010100:	xpb = 256'h0280000002800000000000000000000002800000000000000280000002800000;
		6'b010101:	xpb = 256'h02a0000002a00000000000000000000002a000000000000002a0000002a00000;
		6'b010110:	xpb = 256'h02c0000002c00000000000000000000002c000000000000002c0000002c00000;
		6'b010111:	xpb = 256'h02e0000002e00000000000000000000002e000000000000002e0000002e00000;
		6'b011000:	xpb = 256'h0300000003000000000000000000000003000000000000000300000003000000;
		6'b011001:	xpb = 256'h0320000003200000000000000000000003200000000000000320000003200000;
		6'b011010:	xpb = 256'h0340000003400000000000000000000003400000000000000340000003400000;
		6'b011011:	xpb = 256'h0360000003600000000000000000000003600000000000000360000003600000;
		6'b011100:	xpb = 256'h0380000003800000000000000000000003800000000000000380000003800000;
		6'b011101:	xpb = 256'h03a0000003a00000000000000000000003a000000000000003a0000003a00000;
		6'b011110:	xpb = 256'h03c0000003c00000000000000000000003c000000000000003c0000003c00000;
		6'b011111:	xpb = 256'h03e0000003e00000000000000000000003e000000000000003e0000003e00000;
		6'b100000:	xpb = 256'h0400000004000000000000000000000004000000000000000400000004000000;
		6'b100001:	xpb = 256'h0420000004200000000000000000000004200000000000000420000004200000;
		6'b100010:	xpb = 256'h0440000004400000000000000000000004400000000000000440000004400000;
		6'b100011:	xpb = 256'h0460000004600000000000000000000004600000000000000460000004600000;
		6'b100100:	xpb = 256'h0480000004800000000000000000000004800000000000000480000004800000;
		6'b100101:	xpb = 256'h04a0000004a00000000000000000000004a000000000000004a0000004a00000;
		6'b100110:	xpb = 256'h04c0000004c00000000000000000000004c000000000000004c0000004c00000;
		6'b100111:	xpb = 256'h04e0000004e00000000000000000000004e000000000000004e0000004e00000;
		6'b101000:	xpb = 256'h0500000005000000000000000000000005000000000000000500000005000000;
		6'b101001:	xpb = 256'h0520000005200000000000000000000005200000000000000520000005200000;
		6'b101010:	xpb = 256'h0540000005400000000000000000000005400000000000000540000005400000;
		6'b101011:	xpb = 256'h0560000005600000000000000000000005600000000000000560000005600000;
		6'b101100:	xpb = 256'h0580000005800000000000000000000005800000000000000580000005800000;
		6'b101101:	xpb = 256'h05a0000005a00000000000000000000005a000000000000005a0000005a00000;
		6'b101110:	xpb = 256'h05c0000005c00000000000000000000005c000000000000005c0000005c00000;
		6'b101111:	xpb = 256'h05e0000005e00000000000000000000005e000000000000005e0000005e00000;
		6'b110000:	xpb = 256'h0600000006000000000000000000000006000000000000000600000006000000;
		6'b110001:	xpb = 256'h0620000006200000000000000000000006200000000000000620000006200000;
		6'b110010:	xpb = 256'h0640000006400000000000000000000006400000000000000640000006400000;
		6'b110011:	xpb = 256'h0660000006600000000000000000000006600000000000000660000006600000;
		6'b110100:	xpb = 256'h0680000006800000000000000000000006800000000000000680000006800000;
		6'b110101:	xpb = 256'h06a0000006a00000000000000000000006a000000000000006a0000006a00000;
		6'b110110:	xpb = 256'h06c0000006c00000000000000000000006c000000000000006c0000006c00000;
		6'b110111:	xpb = 256'h06e0000006e00000000000000000000006e000000000000006e0000006e00000;
		6'b111000:	xpb = 256'h0700000007000000000000000000000007000000000000000700000007000000;
		6'b111001:	xpb = 256'h0720000007200000000000000000000007200000000000000720000007200000;
		6'b111010:	xpb = 256'h0740000007400000000000000000000007400000000000000740000007400000;
		6'b111011:	xpb = 256'h0760000007600000000000000000000007600000000000000760000007600000;
		6'b111100:	xpb = 256'h0780000007800000000000000000000007800000000000000780000007800000;
		6'b111101:	xpb = 256'h07a0000007a00000000000000000000007a000000000000007a0000007a00000;
		6'b111110:	xpb = 256'h07c0000007c00000000000000000000007c000000000000007c0000007c00000;
		6'b111111:	xpb = 256'h07e0000007e00000000000000000000007e000000000000007e0000007e00000;
	endcase
end
endmodule

module xpb_23_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0800000008000000000000000000000008000000000000000800000008000000;
		6'b000010:	xpb = 256'h1000000010000000000000000000000010000000000000001000000010000000;
		6'b000011:	xpb = 256'h1800000018000000000000000000000018000000000000001800000018000000;
		6'b000100:	xpb = 256'h2000000020000000000000000000000020000000000000002000000020000000;
		6'b000101:	xpb = 256'h2800000028000000000000000000000028000000000000002800000028000000;
		6'b000110:	xpb = 256'h3000000030000000000000000000000030000000000000003000000030000000;
		6'b000111:	xpb = 256'h3800000038000000000000000000000038000000000000003800000038000000;
		6'b001000:	xpb = 256'h4000000040000000000000000000000040000000000000004000000040000000;
		6'b001001:	xpb = 256'h4800000048000000000000000000000048000000000000004800000048000000;
		6'b001010:	xpb = 256'h5000000050000000000000000000000050000000000000005000000050000000;
		6'b001011:	xpb = 256'h5800000058000000000000000000000058000000000000005800000058000000;
		6'b001100:	xpb = 256'h6000000060000000000000000000000060000000000000006000000060000000;
		6'b001101:	xpb = 256'h6800000068000000000000000000000068000000000000006800000068000000;
		6'b001110:	xpb = 256'h7000000070000000000000000000000070000000000000007000000070000000;
		6'b001111:	xpb = 256'h7800000078000000000000000000000078000000000000007800000078000000;
		6'b010000:	xpb = 256'h8000000080000000000000000000000080000000000000008000000080000000;
		6'b010001:	xpb = 256'h8800000088000000000000000000000088000000000000008800000088000000;
		6'b010010:	xpb = 256'h9000000090000000000000000000000090000000000000009000000090000000;
		6'b010011:	xpb = 256'h9800000098000000000000000000000098000000000000009800000098000000;
		6'b010100:	xpb = 256'ha0000000a00000000000000000000000a000000000000000a0000000a0000000;
		6'b010101:	xpb = 256'ha8000000a80000000000000000000000a800000000000000a8000000a8000000;
		6'b010110:	xpb = 256'hb0000000b00000000000000000000000b000000000000000b0000000b0000000;
		6'b010111:	xpb = 256'hb8000000b80000000000000000000000b800000000000000b8000000b8000000;
		6'b011000:	xpb = 256'hc0000000c00000000000000000000000c000000000000000c0000000c0000000;
		6'b011001:	xpb = 256'hc8000000c80000000000000000000000c800000000000000c8000000c8000000;
		6'b011010:	xpb = 256'hd0000000d00000000000000000000000d000000000000000d0000000d0000000;
		6'b011011:	xpb = 256'hd8000000d80000000000000000000000d800000000000000d8000000d8000000;
		6'b011100:	xpb = 256'he0000000e00000000000000000000000e000000000000000e0000000e0000000;
		6'b011101:	xpb = 256'he8000000e80000000000000000000000e800000000000000e8000000e8000000;
		6'b011110:	xpb = 256'hf0000000f00000000000000000000000f000000000000000f0000000f0000000;
		6'b011111:	xpb = 256'hf8000000f80000000000000000000000f800000000000000f8000000f8000000;
		6'b100000:	xpb = 256'h0000000200000000000000000000000100000001000000000000000100000001;
		6'b100001:	xpb = 256'h0800000208000000000000000000000108000001000000000800000108000001;
		6'b100010:	xpb = 256'h1000000210000000000000000000000110000001000000001000000110000001;
		6'b100011:	xpb = 256'h1800000218000000000000000000000118000001000000001800000118000001;
		6'b100100:	xpb = 256'h2000000220000000000000000000000120000001000000002000000120000001;
		6'b100101:	xpb = 256'h2800000228000000000000000000000128000001000000002800000128000001;
		6'b100110:	xpb = 256'h3000000230000000000000000000000130000001000000003000000130000001;
		6'b100111:	xpb = 256'h3800000238000000000000000000000138000001000000003800000138000001;
		6'b101000:	xpb = 256'h4000000240000000000000000000000140000001000000004000000140000001;
		6'b101001:	xpb = 256'h4800000248000000000000000000000148000001000000004800000148000001;
		6'b101010:	xpb = 256'h5000000250000000000000000000000150000001000000005000000150000001;
		6'b101011:	xpb = 256'h5800000258000000000000000000000158000001000000005800000158000001;
		6'b101100:	xpb = 256'h6000000260000000000000000000000160000001000000006000000160000001;
		6'b101101:	xpb = 256'h6800000268000000000000000000000168000001000000006800000168000001;
		6'b101110:	xpb = 256'h7000000270000000000000000000000170000001000000007000000170000001;
		6'b101111:	xpb = 256'h7800000278000000000000000000000178000001000000007800000178000001;
		6'b110000:	xpb = 256'h8000000280000000000000000000000180000001000000008000000180000001;
		6'b110001:	xpb = 256'h8800000288000000000000000000000188000001000000008800000188000001;
		6'b110010:	xpb = 256'h9000000290000000000000000000000190000001000000009000000190000001;
		6'b110011:	xpb = 256'h9800000298000000000000000000000198000001000000009800000198000001;
		6'b110100:	xpb = 256'ha0000002a00000000000000000000001a000000100000000a0000001a0000001;
		6'b110101:	xpb = 256'ha8000002a80000000000000000000001a800000100000000a8000001a8000001;
		6'b110110:	xpb = 256'hb0000002b00000000000000000000001b000000100000000b0000001b0000001;
		6'b110111:	xpb = 256'hb8000002b80000000000000000000001b800000100000000b8000001b8000001;
		6'b111000:	xpb = 256'hc0000002c00000000000000000000001c000000100000000c0000001c0000001;
		6'b111001:	xpb = 256'hc8000002c80000000000000000000001c800000100000000c8000001c8000001;
		6'b111010:	xpb = 256'hd0000002d00000000000000000000001d000000100000000d0000001d0000001;
		6'b111011:	xpb = 256'hd8000002d80000000000000000000001d800000100000000d8000001d8000001;
		6'b111100:	xpb = 256'he0000002e00000000000000000000001e000000100000000e0000001e0000001;
		6'b111101:	xpb = 256'he8000002e80000000000000000000001e800000100000000e8000001e8000001;
		6'b111110:	xpb = 256'hf0000002f00000000000000000000001f000000100000000f0000001f0000001;
		6'b111111:	xpb = 256'hf8000002f80000000000000000000001f800000100000000f8000001f8000001;
	endcase
end
endmodule

module xpb_24_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000200000000000000000000000100000001000000000000000100000001;
		5'b00010:	xpb = 256'h0000000400000000000000000000000200000002000000000000000200000002;
		5'b00011:	xpb = 256'h0000000600000000000000000000000300000003000000000000000300000003;
		5'b00100:	xpb = 256'h0000000800000000000000000000000400000004000000000000000400000004;
		5'b00101:	xpb = 256'h0000000a00000000000000000000000500000005000000000000000500000005;
		5'b00110:	xpb = 256'h0000000c00000000000000000000000600000006000000000000000600000006;
		5'b00111:	xpb = 256'h0000000e00000000000000000000000700000007000000000000000700000007;
		5'b01000:	xpb = 256'h0000001000000000000000000000000800000008000000000000000800000008;
		5'b01001:	xpb = 256'h0000001200000000000000000000000900000009000000000000000900000009;
		5'b01010:	xpb = 256'h0000001400000000000000000000000a0000000a000000000000000a0000000a;
		5'b01011:	xpb = 256'h0000001600000000000000000000000b0000000b000000000000000b0000000b;
		5'b01100:	xpb = 256'h0000001800000000000000000000000c0000000c000000000000000c0000000c;
		5'b01101:	xpb = 256'h0000001a00000000000000000000000d0000000d000000000000000d0000000d;
		5'b01110:	xpb = 256'h0000001c00000000000000000000000e0000000e000000000000000e0000000e;
		5'b01111:	xpb = 256'h0000001e00000000000000000000000f0000000f000000000000000f0000000f;
		5'b10000:	xpb = 256'h0000002000000000000000000000001000000010000000000000001000000010;
		5'b10001:	xpb = 256'h0000002200000000000000000000001100000011000000000000001100000011;
		5'b10010:	xpb = 256'h0000002400000000000000000000001200000012000000000000001200000012;
		5'b10011:	xpb = 256'h0000002600000000000000000000001300000013000000000000001300000013;
		5'b10100:	xpb = 256'h0000002800000000000000000000001400000014000000000000001400000014;
		5'b10101:	xpb = 256'h0000002a00000000000000000000001500000015000000000000001500000015;
		5'b10110:	xpb = 256'h0000002c00000000000000000000001600000016000000000000001600000016;
		5'b10111:	xpb = 256'h0000002e00000000000000000000001700000017000000000000001700000017;
		5'b11000:	xpb = 256'h0000003000000000000000000000001800000018000000000000001800000018;
		5'b11001:	xpb = 256'h0000003200000000000000000000001900000019000000000000001900000019;
		5'b11010:	xpb = 256'h0000003400000000000000000000001a0000001a000000000000001a0000001a;
		5'b11011:	xpb = 256'h0000003600000000000000000000001b0000001b000000000000001b0000001b;
		5'b11100:	xpb = 256'h0000003800000000000000000000001c0000001c000000000000001c0000001c;
		5'b11101:	xpb = 256'h0000003a00000000000000000000001d0000001d000000000000001d0000001d;
		5'b11110:	xpb = 256'h0000003c00000000000000000000001e0000001e000000000000001e0000001e;
		5'b11111:	xpb = 256'h0000003e00000000000000000000001f0000001f000000000000001f0000001f;
	endcase
end
endmodule

module xpb_24_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000004000000000000000000000002000000020000000000000002000000020;
		6'b000010:	xpb = 256'h0000008000000000000000000000004000000040000000000000004000000040;
		6'b000011:	xpb = 256'h000000c000000000000000000000006000000060000000000000006000000060;
		6'b000100:	xpb = 256'h0000010000000000000000000000008000000080000000000000008000000080;
		6'b000101:	xpb = 256'h000001400000000000000000000000a0000000a000000000000000a0000000a0;
		6'b000110:	xpb = 256'h000001800000000000000000000000c0000000c000000000000000c0000000c0;
		6'b000111:	xpb = 256'h000001c00000000000000000000000e0000000e000000000000000e0000000e0;
		6'b001000:	xpb = 256'h0000020000000000000000000000010000000100000000000000010000000100;
		6'b001001:	xpb = 256'h0000024000000000000000000000012000000120000000000000012000000120;
		6'b001010:	xpb = 256'h0000028000000000000000000000014000000140000000000000014000000140;
		6'b001011:	xpb = 256'h000002c000000000000000000000016000000160000000000000016000000160;
		6'b001100:	xpb = 256'h0000030000000000000000000000018000000180000000000000018000000180;
		6'b001101:	xpb = 256'h000003400000000000000000000001a0000001a000000000000001a0000001a0;
		6'b001110:	xpb = 256'h000003800000000000000000000001c0000001c000000000000001c0000001c0;
		6'b001111:	xpb = 256'h000003c00000000000000000000001e0000001e000000000000001e0000001e0;
		6'b010000:	xpb = 256'h0000040000000000000000000000020000000200000000000000020000000200;
		6'b010001:	xpb = 256'h0000044000000000000000000000022000000220000000000000022000000220;
		6'b010010:	xpb = 256'h0000048000000000000000000000024000000240000000000000024000000240;
		6'b010011:	xpb = 256'h000004c000000000000000000000026000000260000000000000026000000260;
		6'b010100:	xpb = 256'h0000050000000000000000000000028000000280000000000000028000000280;
		6'b010101:	xpb = 256'h000005400000000000000000000002a0000002a000000000000002a0000002a0;
		6'b010110:	xpb = 256'h000005800000000000000000000002c0000002c000000000000002c0000002c0;
		6'b010111:	xpb = 256'h000005c00000000000000000000002e0000002e000000000000002e0000002e0;
		6'b011000:	xpb = 256'h0000060000000000000000000000030000000300000000000000030000000300;
		6'b011001:	xpb = 256'h0000064000000000000000000000032000000320000000000000032000000320;
		6'b011010:	xpb = 256'h0000068000000000000000000000034000000340000000000000034000000340;
		6'b011011:	xpb = 256'h000006c000000000000000000000036000000360000000000000036000000360;
		6'b011100:	xpb = 256'h0000070000000000000000000000038000000380000000000000038000000380;
		6'b011101:	xpb = 256'h000007400000000000000000000003a0000003a000000000000003a0000003a0;
		6'b011110:	xpb = 256'h000007800000000000000000000003c0000003c000000000000003c0000003c0;
		6'b011111:	xpb = 256'h000007c00000000000000000000003e0000003e000000000000003e0000003e0;
		6'b100000:	xpb = 256'h0000080000000000000000000000040000000400000000000000040000000400;
		6'b100001:	xpb = 256'h0000084000000000000000000000042000000420000000000000042000000420;
		6'b100010:	xpb = 256'h0000088000000000000000000000044000000440000000000000044000000440;
		6'b100011:	xpb = 256'h000008c000000000000000000000046000000460000000000000046000000460;
		6'b100100:	xpb = 256'h0000090000000000000000000000048000000480000000000000048000000480;
		6'b100101:	xpb = 256'h000009400000000000000000000004a0000004a000000000000004a0000004a0;
		6'b100110:	xpb = 256'h000009800000000000000000000004c0000004c000000000000004c0000004c0;
		6'b100111:	xpb = 256'h000009c00000000000000000000004e0000004e000000000000004e0000004e0;
		6'b101000:	xpb = 256'h00000a0000000000000000000000050000000500000000000000050000000500;
		6'b101001:	xpb = 256'h00000a4000000000000000000000052000000520000000000000052000000520;
		6'b101010:	xpb = 256'h00000a8000000000000000000000054000000540000000000000054000000540;
		6'b101011:	xpb = 256'h00000ac000000000000000000000056000000560000000000000056000000560;
		6'b101100:	xpb = 256'h00000b0000000000000000000000058000000580000000000000058000000580;
		6'b101101:	xpb = 256'h00000b400000000000000000000005a0000005a000000000000005a0000005a0;
		6'b101110:	xpb = 256'h00000b800000000000000000000005c0000005c000000000000005c0000005c0;
		6'b101111:	xpb = 256'h00000bc00000000000000000000005e0000005e000000000000005e0000005e0;
		6'b110000:	xpb = 256'h00000c0000000000000000000000060000000600000000000000060000000600;
		6'b110001:	xpb = 256'h00000c4000000000000000000000062000000620000000000000062000000620;
		6'b110010:	xpb = 256'h00000c8000000000000000000000064000000640000000000000064000000640;
		6'b110011:	xpb = 256'h00000cc000000000000000000000066000000660000000000000066000000660;
		6'b110100:	xpb = 256'h00000d0000000000000000000000068000000680000000000000068000000680;
		6'b110101:	xpb = 256'h00000d400000000000000000000006a0000006a000000000000006a0000006a0;
		6'b110110:	xpb = 256'h00000d800000000000000000000006c0000006c000000000000006c0000006c0;
		6'b110111:	xpb = 256'h00000dc00000000000000000000006e0000006e000000000000006e0000006e0;
		6'b111000:	xpb = 256'h00000e0000000000000000000000070000000700000000000000070000000700;
		6'b111001:	xpb = 256'h00000e4000000000000000000000072000000720000000000000072000000720;
		6'b111010:	xpb = 256'h00000e8000000000000000000000074000000740000000000000074000000740;
		6'b111011:	xpb = 256'h00000ec000000000000000000000076000000760000000000000076000000760;
		6'b111100:	xpb = 256'h00000f0000000000000000000000078000000780000000000000078000000780;
		6'b111101:	xpb = 256'h00000f400000000000000000000007a0000007a000000000000007a0000007a0;
		6'b111110:	xpb = 256'h00000f800000000000000000000007c0000007c000000000000007c0000007c0;
		6'b111111:	xpb = 256'h00000fc00000000000000000000007e0000007e000000000000007e0000007e0;
	endcase
end
endmodule

module xpb_24_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000100000000000000000000000080000000800000000000000080000000800;
		6'b000010:	xpb = 256'h0000200000000000000000000000100000001000000000000000100000001000;
		6'b000011:	xpb = 256'h0000300000000000000000000000180000001800000000000000180000001800;
		6'b000100:	xpb = 256'h0000400000000000000000000000200000002000000000000000200000002000;
		6'b000101:	xpb = 256'h0000500000000000000000000000280000002800000000000000280000002800;
		6'b000110:	xpb = 256'h0000600000000000000000000000300000003000000000000000300000003000;
		6'b000111:	xpb = 256'h0000700000000000000000000000380000003800000000000000380000003800;
		6'b001000:	xpb = 256'h0000800000000000000000000000400000004000000000000000400000004000;
		6'b001001:	xpb = 256'h0000900000000000000000000000480000004800000000000000480000004800;
		6'b001010:	xpb = 256'h0000a00000000000000000000000500000005000000000000000500000005000;
		6'b001011:	xpb = 256'h0000b00000000000000000000000580000005800000000000000580000005800;
		6'b001100:	xpb = 256'h0000c00000000000000000000000600000006000000000000000600000006000;
		6'b001101:	xpb = 256'h0000d00000000000000000000000680000006800000000000000680000006800;
		6'b001110:	xpb = 256'h0000e00000000000000000000000700000007000000000000000700000007000;
		6'b001111:	xpb = 256'h0000f00000000000000000000000780000007800000000000000780000007800;
		6'b010000:	xpb = 256'h0001000000000000000000000000800000008000000000000000800000008000;
		6'b010001:	xpb = 256'h0001100000000000000000000000880000008800000000000000880000008800;
		6'b010010:	xpb = 256'h0001200000000000000000000000900000009000000000000000900000009000;
		6'b010011:	xpb = 256'h0001300000000000000000000000980000009800000000000000980000009800;
		6'b010100:	xpb = 256'h0001400000000000000000000000a0000000a000000000000000a0000000a000;
		6'b010101:	xpb = 256'h0001500000000000000000000000a8000000a800000000000000a8000000a800;
		6'b010110:	xpb = 256'h0001600000000000000000000000b0000000b000000000000000b0000000b000;
		6'b010111:	xpb = 256'h0001700000000000000000000000b8000000b800000000000000b8000000b800;
		6'b011000:	xpb = 256'h0001800000000000000000000000c0000000c000000000000000c0000000c000;
		6'b011001:	xpb = 256'h0001900000000000000000000000c8000000c800000000000000c8000000c800;
		6'b011010:	xpb = 256'h0001a00000000000000000000000d0000000d000000000000000d0000000d000;
		6'b011011:	xpb = 256'h0001b00000000000000000000000d8000000d800000000000000d8000000d800;
		6'b011100:	xpb = 256'h0001c00000000000000000000000e0000000e000000000000000e0000000e000;
		6'b011101:	xpb = 256'h0001d00000000000000000000000e8000000e800000000000000e8000000e800;
		6'b011110:	xpb = 256'h0001e00000000000000000000000f0000000f000000000000000f0000000f000;
		6'b011111:	xpb = 256'h0001f00000000000000000000000f8000000f800000000000000f8000000f800;
		6'b100000:	xpb = 256'h0002000000000000000000000001000000010000000000000001000000010000;
		6'b100001:	xpb = 256'h0002100000000000000000000001080000010800000000000001080000010800;
		6'b100010:	xpb = 256'h0002200000000000000000000001100000011000000000000001100000011000;
		6'b100011:	xpb = 256'h0002300000000000000000000001180000011800000000000001180000011800;
		6'b100100:	xpb = 256'h0002400000000000000000000001200000012000000000000001200000012000;
		6'b100101:	xpb = 256'h0002500000000000000000000001280000012800000000000001280000012800;
		6'b100110:	xpb = 256'h0002600000000000000000000001300000013000000000000001300000013000;
		6'b100111:	xpb = 256'h0002700000000000000000000001380000013800000000000001380000013800;
		6'b101000:	xpb = 256'h0002800000000000000000000001400000014000000000000001400000014000;
		6'b101001:	xpb = 256'h0002900000000000000000000001480000014800000000000001480000014800;
		6'b101010:	xpb = 256'h0002a00000000000000000000001500000015000000000000001500000015000;
		6'b101011:	xpb = 256'h0002b00000000000000000000001580000015800000000000001580000015800;
		6'b101100:	xpb = 256'h0002c00000000000000000000001600000016000000000000001600000016000;
		6'b101101:	xpb = 256'h0002d00000000000000000000001680000016800000000000001680000016800;
		6'b101110:	xpb = 256'h0002e00000000000000000000001700000017000000000000001700000017000;
		6'b101111:	xpb = 256'h0002f00000000000000000000001780000017800000000000001780000017800;
		6'b110000:	xpb = 256'h0003000000000000000000000001800000018000000000000001800000018000;
		6'b110001:	xpb = 256'h0003100000000000000000000001880000018800000000000001880000018800;
		6'b110010:	xpb = 256'h0003200000000000000000000001900000019000000000000001900000019000;
		6'b110011:	xpb = 256'h0003300000000000000000000001980000019800000000000001980000019800;
		6'b110100:	xpb = 256'h0003400000000000000000000001a0000001a000000000000001a0000001a000;
		6'b110101:	xpb = 256'h0003500000000000000000000001a8000001a800000000000001a8000001a800;
		6'b110110:	xpb = 256'h0003600000000000000000000001b0000001b000000000000001b0000001b000;
		6'b110111:	xpb = 256'h0003700000000000000000000001b8000001b800000000000001b8000001b800;
		6'b111000:	xpb = 256'h0003800000000000000000000001c0000001c000000000000001c0000001c000;
		6'b111001:	xpb = 256'h0003900000000000000000000001c8000001c800000000000001c8000001c800;
		6'b111010:	xpb = 256'h0003a00000000000000000000001d0000001d000000000000001d0000001d000;
		6'b111011:	xpb = 256'h0003b00000000000000000000001d8000001d800000000000001d8000001d800;
		6'b111100:	xpb = 256'h0003c00000000000000000000001e0000001e000000000000001e0000001e000;
		6'b111101:	xpb = 256'h0003d00000000000000000000001e8000001e800000000000001e8000001e800;
		6'b111110:	xpb = 256'h0003e00000000000000000000001f0000001f000000000000001f0000001f000;
		6'b111111:	xpb = 256'h0003f00000000000000000000001f8000001f800000000000001f8000001f800;
	endcase
end
endmodule

module xpb_25_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0002000000000000000000000001000000010000000000000001000000010000;
		5'b00010:	xpb = 256'h0004000000000000000000000002000000020000000000000002000000020000;
		5'b00011:	xpb = 256'h0006000000000000000000000003000000030000000000000003000000030000;
		5'b00100:	xpb = 256'h0008000000000000000000000004000000040000000000000004000000040000;
		5'b00101:	xpb = 256'h000a000000000000000000000005000000050000000000000005000000050000;
		5'b00110:	xpb = 256'h000c000000000000000000000006000000060000000000000006000000060000;
		5'b00111:	xpb = 256'h000e000000000000000000000007000000070000000000000007000000070000;
		5'b01000:	xpb = 256'h0010000000000000000000000008000000080000000000000008000000080000;
		5'b01001:	xpb = 256'h0012000000000000000000000009000000090000000000000009000000090000;
		5'b01010:	xpb = 256'h001400000000000000000000000a0000000a000000000000000a0000000a0000;
		5'b01011:	xpb = 256'h001600000000000000000000000b0000000b000000000000000b0000000b0000;
		5'b01100:	xpb = 256'h001800000000000000000000000c0000000c000000000000000c0000000c0000;
		5'b01101:	xpb = 256'h001a00000000000000000000000d0000000d000000000000000d0000000d0000;
		5'b01110:	xpb = 256'h001c00000000000000000000000e0000000e000000000000000e0000000e0000;
		5'b01111:	xpb = 256'h001e00000000000000000000000f0000000f000000000000000f0000000f0000;
		5'b10000:	xpb = 256'h0020000000000000000000000010000000100000000000000010000000100000;
		5'b10001:	xpb = 256'h0022000000000000000000000011000000110000000000000011000000110000;
		5'b10010:	xpb = 256'h0024000000000000000000000012000000120000000000000012000000120000;
		5'b10011:	xpb = 256'h0026000000000000000000000013000000130000000000000013000000130000;
		5'b10100:	xpb = 256'h0028000000000000000000000014000000140000000000000014000000140000;
		5'b10101:	xpb = 256'h002a000000000000000000000015000000150000000000000015000000150000;
		5'b10110:	xpb = 256'h002c000000000000000000000016000000160000000000000016000000160000;
		5'b10111:	xpb = 256'h002e000000000000000000000017000000170000000000000017000000170000;
		5'b11000:	xpb = 256'h0030000000000000000000000018000000180000000000000018000000180000;
		5'b11001:	xpb = 256'h0032000000000000000000000019000000190000000000000019000000190000;
		5'b11010:	xpb = 256'h003400000000000000000000001a0000001a000000000000001a0000001a0000;
		5'b11011:	xpb = 256'h003600000000000000000000001b0000001b000000000000001b0000001b0000;
		5'b11100:	xpb = 256'h003800000000000000000000001c0000001c000000000000001c0000001c0000;
		5'b11101:	xpb = 256'h003a00000000000000000000001d0000001d000000000000001d0000001d0000;
		5'b11110:	xpb = 256'h003c00000000000000000000001e0000001e000000000000001e0000001e0000;
		5'b11111:	xpb = 256'h003e00000000000000000000001f0000001f000000000000001f0000001f0000;
	endcase
end
endmodule

module xpb_25_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0040000000000000000000000020000000200000000000000020000000200000;
		6'b000010:	xpb = 256'h0080000000000000000000000040000000400000000000000040000000400000;
		6'b000011:	xpb = 256'h00c0000000000000000000000060000000600000000000000060000000600000;
		6'b000100:	xpb = 256'h0100000000000000000000000080000000800000000000000080000000800000;
		6'b000101:	xpb = 256'h01400000000000000000000000a0000000a000000000000000a0000000a00000;
		6'b000110:	xpb = 256'h01800000000000000000000000c0000000c000000000000000c0000000c00000;
		6'b000111:	xpb = 256'h01c00000000000000000000000e0000000e000000000000000e0000000e00000;
		6'b001000:	xpb = 256'h0200000000000000000000000100000001000000000000000100000001000000;
		6'b001001:	xpb = 256'h0240000000000000000000000120000001200000000000000120000001200000;
		6'b001010:	xpb = 256'h0280000000000000000000000140000001400000000000000140000001400000;
		6'b001011:	xpb = 256'h02c0000000000000000000000160000001600000000000000160000001600000;
		6'b001100:	xpb = 256'h0300000000000000000000000180000001800000000000000180000001800000;
		6'b001101:	xpb = 256'h03400000000000000000000001a0000001a000000000000001a0000001a00000;
		6'b001110:	xpb = 256'h03800000000000000000000001c0000001c000000000000001c0000001c00000;
		6'b001111:	xpb = 256'h03c00000000000000000000001e0000001e000000000000001e0000001e00000;
		6'b010000:	xpb = 256'h0400000000000000000000000200000002000000000000000200000002000000;
		6'b010001:	xpb = 256'h0440000000000000000000000220000002200000000000000220000002200000;
		6'b010010:	xpb = 256'h0480000000000000000000000240000002400000000000000240000002400000;
		6'b010011:	xpb = 256'h04c0000000000000000000000260000002600000000000000260000002600000;
		6'b010100:	xpb = 256'h0500000000000000000000000280000002800000000000000280000002800000;
		6'b010101:	xpb = 256'h05400000000000000000000002a0000002a000000000000002a0000002a00000;
		6'b010110:	xpb = 256'h05800000000000000000000002c0000002c000000000000002c0000002c00000;
		6'b010111:	xpb = 256'h05c00000000000000000000002e0000002e000000000000002e0000002e00000;
		6'b011000:	xpb = 256'h0600000000000000000000000300000003000000000000000300000003000000;
		6'b011001:	xpb = 256'h0640000000000000000000000320000003200000000000000320000003200000;
		6'b011010:	xpb = 256'h0680000000000000000000000340000003400000000000000340000003400000;
		6'b011011:	xpb = 256'h06c0000000000000000000000360000003600000000000000360000003600000;
		6'b011100:	xpb = 256'h0700000000000000000000000380000003800000000000000380000003800000;
		6'b011101:	xpb = 256'h07400000000000000000000003a0000003a000000000000003a0000003a00000;
		6'b011110:	xpb = 256'h07800000000000000000000003c0000003c000000000000003c0000003c00000;
		6'b011111:	xpb = 256'h07c00000000000000000000003e0000003e000000000000003e0000003e00000;
		6'b100000:	xpb = 256'h0800000000000000000000000400000004000000000000000400000004000000;
		6'b100001:	xpb = 256'h0840000000000000000000000420000004200000000000000420000004200000;
		6'b100010:	xpb = 256'h0880000000000000000000000440000004400000000000000440000004400000;
		6'b100011:	xpb = 256'h08c0000000000000000000000460000004600000000000000460000004600000;
		6'b100100:	xpb = 256'h0900000000000000000000000480000004800000000000000480000004800000;
		6'b100101:	xpb = 256'h09400000000000000000000004a0000004a000000000000004a0000004a00000;
		6'b100110:	xpb = 256'h09800000000000000000000004c0000004c000000000000004c0000004c00000;
		6'b100111:	xpb = 256'h09c00000000000000000000004e0000004e000000000000004e0000004e00000;
		6'b101000:	xpb = 256'h0a00000000000000000000000500000005000000000000000500000005000000;
		6'b101001:	xpb = 256'h0a40000000000000000000000520000005200000000000000520000005200000;
		6'b101010:	xpb = 256'h0a80000000000000000000000540000005400000000000000540000005400000;
		6'b101011:	xpb = 256'h0ac0000000000000000000000560000005600000000000000560000005600000;
		6'b101100:	xpb = 256'h0b00000000000000000000000580000005800000000000000580000005800000;
		6'b101101:	xpb = 256'h0b400000000000000000000005a0000005a000000000000005a0000005a00000;
		6'b101110:	xpb = 256'h0b800000000000000000000005c0000005c000000000000005c0000005c00000;
		6'b101111:	xpb = 256'h0bc00000000000000000000005e0000005e000000000000005e0000005e00000;
		6'b110000:	xpb = 256'h0c00000000000000000000000600000006000000000000000600000006000000;
		6'b110001:	xpb = 256'h0c40000000000000000000000620000006200000000000000620000006200000;
		6'b110010:	xpb = 256'h0c80000000000000000000000640000006400000000000000640000006400000;
		6'b110011:	xpb = 256'h0cc0000000000000000000000660000006600000000000000660000006600000;
		6'b110100:	xpb = 256'h0d00000000000000000000000680000006800000000000000680000006800000;
		6'b110101:	xpb = 256'h0d400000000000000000000006a0000006a000000000000006a0000006a00000;
		6'b110110:	xpb = 256'h0d800000000000000000000006c0000006c000000000000006c0000006c00000;
		6'b110111:	xpb = 256'h0dc00000000000000000000006e0000006e000000000000006e0000006e00000;
		6'b111000:	xpb = 256'h0e00000000000000000000000700000007000000000000000700000007000000;
		6'b111001:	xpb = 256'h0e40000000000000000000000720000007200000000000000720000007200000;
		6'b111010:	xpb = 256'h0e80000000000000000000000740000007400000000000000740000007400000;
		6'b111011:	xpb = 256'h0ec0000000000000000000000760000007600000000000000760000007600000;
		6'b111100:	xpb = 256'h0f00000000000000000000000780000007800000000000000780000007800000;
		6'b111101:	xpb = 256'h0f400000000000000000000007a0000007a000000000000007a0000007a00000;
		6'b111110:	xpb = 256'h0f800000000000000000000007c0000007c000000000000007c0000007c00000;
		6'b111111:	xpb = 256'h0fc00000000000000000000007e0000007e000000000000007e0000007e00000;
	endcase
end
endmodule

module xpb_25_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h1000000000000000000000000800000008000000000000000800000008000000;
		6'b000010:	xpb = 256'h2000000000000000000000001000000010000000000000001000000010000000;
		6'b000011:	xpb = 256'h3000000000000000000000001800000018000000000000001800000018000000;
		6'b000100:	xpb = 256'h4000000000000000000000002000000020000000000000002000000020000000;
		6'b000101:	xpb = 256'h5000000000000000000000002800000028000000000000002800000028000000;
		6'b000110:	xpb = 256'h6000000000000000000000003000000030000000000000003000000030000000;
		6'b000111:	xpb = 256'h7000000000000000000000003800000038000000000000003800000038000000;
		6'b001000:	xpb = 256'h8000000000000000000000004000000040000000000000004000000040000000;
		6'b001001:	xpb = 256'h9000000000000000000000004800000048000000000000004800000048000000;
		6'b001010:	xpb = 256'ha000000000000000000000005000000050000000000000005000000050000000;
		6'b001011:	xpb = 256'hb000000000000000000000005800000058000000000000005800000058000000;
		6'b001100:	xpb = 256'hc000000000000000000000006000000060000000000000006000000060000000;
		6'b001101:	xpb = 256'hd000000000000000000000006800000068000000000000006800000068000000;
		6'b001110:	xpb = 256'he000000000000000000000007000000070000000000000007000000070000000;
		6'b001111:	xpb = 256'hf000000000000000000000007800000078000000000000007800000078000000;
		6'b010000:	xpb = 256'h0000000100000000000000008000000080000000ffffffff8000000080000001;
		6'b010001:	xpb = 256'h1000000100000000000000008800000088000000ffffffff8800000088000001;
		6'b010010:	xpb = 256'h2000000100000000000000009000000090000000ffffffff9000000090000001;
		6'b010011:	xpb = 256'h3000000100000000000000009800000098000000ffffffff9800000098000001;
		6'b010100:	xpb = 256'h400000010000000000000000a0000000a0000000ffffffffa0000000a0000001;
		6'b010101:	xpb = 256'h500000010000000000000000a8000000a8000000ffffffffa8000000a8000001;
		6'b010110:	xpb = 256'h600000010000000000000000b0000000b0000000ffffffffb0000000b0000001;
		6'b010111:	xpb = 256'h700000010000000000000000b8000000b8000000ffffffffb8000000b8000001;
		6'b011000:	xpb = 256'h800000010000000000000000c0000000c0000000ffffffffc0000000c0000001;
		6'b011001:	xpb = 256'h900000010000000000000000c8000000c8000000ffffffffc8000000c8000001;
		6'b011010:	xpb = 256'ha00000010000000000000000d0000000d0000000ffffffffd0000000d0000001;
		6'b011011:	xpb = 256'hb00000010000000000000000d8000000d8000000ffffffffd8000000d8000001;
		6'b011100:	xpb = 256'hc00000010000000000000000e0000000e0000000ffffffffe0000000e0000001;
		6'b011101:	xpb = 256'hd00000010000000000000000e8000000e8000000ffffffffe8000000e8000001;
		6'b011110:	xpb = 256'he00000010000000000000000f0000000f0000000fffffffff0000000f0000001;
		6'b011111:	xpb = 256'hf00000010000000000000000f8000000f8000000fffffffff8000000f8000001;
		6'b100000:	xpb = 256'h0000000200000000000000010000000100000001ffffffff0000000100000002;
		6'b100001:	xpb = 256'h1000000200000000000000010800000108000001ffffffff0800000108000002;
		6'b100010:	xpb = 256'h2000000200000000000000011000000110000001ffffffff1000000110000002;
		6'b100011:	xpb = 256'h3000000200000000000000011800000118000001ffffffff1800000118000002;
		6'b100100:	xpb = 256'h4000000200000000000000012000000120000001ffffffff2000000120000002;
		6'b100101:	xpb = 256'h5000000200000000000000012800000128000001ffffffff2800000128000002;
		6'b100110:	xpb = 256'h6000000200000000000000013000000130000001ffffffff3000000130000002;
		6'b100111:	xpb = 256'h7000000200000000000000013800000138000001ffffffff3800000138000002;
		6'b101000:	xpb = 256'h8000000200000000000000014000000140000001ffffffff4000000140000002;
		6'b101001:	xpb = 256'h9000000200000000000000014800000148000001ffffffff4800000148000002;
		6'b101010:	xpb = 256'ha000000200000000000000015000000150000001ffffffff5000000150000002;
		6'b101011:	xpb = 256'hb000000200000000000000015800000158000001ffffffff5800000158000002;
		6'b101100:	xpb = 256'hc000000200000000000000016000000160000001ffffffff6000000160000002;
		6'b101101:	xpb = 256'hd000000200000000000000016800000168000001ffffffff6800000168000002;
		6'b101110:	xpb = 256'he000000200000000000000017000000170000001ffffffff7000000170000002;
		6'b101111:	xpb = 256'hf000000200000000000000017800000178000001ffffffff7800000178000002;
		6'b110000:	xpb = 256'h0000000300000000000000018000000180000002fffffffe8000000180000003;
		6'b110001:	xpb = 256'h1000000300000000000000018800000188000002fffffffe8800000188000003;
		6'b110010:	xpb = 256'h2000000300000000000000019000000190000002fffffffe9000000190000003;
		6'b110011:	xpb = 256'h3000000300000000000000019800000198000002fffffffe9800000198000003;
		6'b110100:	xpb = 256'h400000030000000000000001a0000001a0000002fffffffea0000001a0000003;
		6'b110101:	xpb = 256'h500000030000000000000001a8000001a8000002fffffffea8000001a8000003;
		6'b110110:	xpb = 256'h600000030000000000000001b0000001b0000002fffffffeb0000001b0000003;
		6'b110111:	xpb = 256'h700000030000000000000001b8000001b8000002fffffffeb8000001b8000003;
		6'b111000:	xpb = 256'h800000030000000000000001c0000001c0000002fffffffec0000001c0000003;
		6'b111001:	xpb = 256'h900000030000000000000001c8000001c8000002fffffffec8000001c8000003;
		6'b111010:	xpb = 256'ha00000030000000000000001d0000001d0000002fffffffed0000001d0000003;
		6'b111011:	xpb = 256'hb00000030000000000000001d8000001d8000002fffffffed8000001d8000003;
		6'b111100:	xpb = 256'hc00000030000000000000001e0000001e0000002fffffffee0000001e0000003;
		6'b111101:	xpb = 256'hd00000030000000000000001e8000001e8000002fffffffee8000001e8000003;
		6'b111110:	xpb = 256'he00000030000000000000001f0000001f0000002fffffffef0000001f0000003;
		6'b111111:	xpb = 256'hf00000030000000000000001f8000001f8000002fffffffef8000001f8000003;
	endcase
end
endmodule

module xpb_26_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000200000000000000010000000100000001ffffffff0000000100000002;
		5'b00010:	xpb = 256'h0000000400000000000000020000000200000003fffffffe0000000200000004;
		5'b00011:	xpb = 256'h0000000600000000000000030000000300000005fffffffd0000000300000006;
		5'b00100:	xpb = 256'h0000000800000000000000040000000400000007fffffffc0000000400000008;
		5'b00101:	xpb = 256'h0000000a00000000000000050000000500000009fffffffb000000050000000a;
		5'b00110:	xpb = 256'h0000000c0000000000000006000000060000000bfffffffa000000060000000c;
		5'b00111:	xpb = 256'h0000000e0000000000000007000000070000000dfffffff9000000070000000e;
		5'b01000:	xpb = 256'h000000100000000000000008000000080000000ffffffff80000000800000010;
		5'b01001:	xpb = 256'h0000001200000000000000090000000900000011fffffff70000000900000012;
		5'b01010:	xpb = 256'h00000014000000000000000a0000000a00000013fffffff60000000a00000014;
		5'b01011:	xpb = 256'h00000016000000000000000b0000000b00000015fffffff50000000b00000016;
		5'b01100:	xpb = 256'h00000018000000000000000c0000000c00000017fffffff40000000c00000018;
		5'b01101:	xpb = 256'h0000001a000000000000000d0000000d00000019fffffff30000000d0000001a;
		5'b01110:	xpb = 256'h0000001c000000000000000e0000000e0000001bfffffff20000000e0000001c;
		5'b01111:	xpb = 256'h0000001e000000000000000f0000000f0000001dfffffff10000000f0000001e;
		5'b10000:	xpb = 256'h000000200000000000000010000000100000001ffffffff00000001000000020;
		5'b10001:	xpb = 256'h0000002200000000000000110000001100000021ffffffef0000001100000022;
		5'b10010:	xpb = 256'h0000002400000000000000120000001200000023ffffffee0000001200000024;
		5'b10011:	xpb = 256'h0000002600000000000000130000001300000025ffffffed0000001300000026;
		5'b10100:	xpb = 256'h0000002800000000000000140000001400000027ffffffec0000001400000028;
		5'b10101:	xpb = 256'h0000002a00000000000000150000001500000029ffffffeb000000150000002a;
		5'b10110:	xpb = 256'h0000002c0000000000000016000000160000002bffffffea000000160000002c;
		5'b10111:	xpb = 256'h0000002e0000000000000017000000170000002dffffffe9000000170000002e;
		5'b11000:	xpb = 256'h000000300000000000000018000000180000002fffffffe80000001800000030;
		5'b11001:	xpb = 256'h0000003200000000000000190000001900000031ffffffe70000001900000032;
		5'b11010:	xpb = 256'h00000034000000000000001a0000001a00000033ffffffe60000001a00000034;
		5'b11011:	xpb = 256'h00000036000000000000001b0000001b00000035ffffffe50000001b00000036;
		5'b11100:	xpb = 256'h00000038000000000000001c0000001c00000037ffffffe40000001c00000038;
		5'b11101:	xpb = 256'h0000003a000000000000001d0000001d00000039ffffffe30000001d0000003a;
		5'b11110:	xpb = 256'h0000003c000000000000001e0000001e0000003bffffffe20000001e0000003c;
		5'b11111:	xpb = 256'h0000003e000000000000001f0000001f0000003dffffffe10000001f0000003e;
	endcase
end
endmodule

module xpb_26_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h000000400000000000000020000000200000003fffffffe00000002000000040;
		6'b000010:	xpb = 256'h000000800000000000000040000000400000007fffffffc00000004000000080;
		6'b000011:	xpb = 256'h000000c0000000000000006000000060000000bfffffffa000000060000000c0;
		6'b000100:	xpb = 256'h00000100000000000000008000000080000000ffffffff800000008000000100;
		6'b000101:	xpb = 256'h0000014000000000000000a0000000a00000013fffffff60000000a000000140;
		6'b000110:	xpb = 256'h0000018000000000000000c0000000c00000017fffffff40000000c000000180;
		6'b000111:	xpb = 256'h000001c000000000000000e0000000e0000001bfffffff20000000e0000001c0;
		6'b001000:	xpb = 256'h00000200000000000000010000000100000001ffffffff000000010000000200;
		6'b001001:	xpb = 256'h000002400000000000000120000001200000023ffffffee00000012000000240;
		6'b001010:	xpb = 256'h000002800000000000000140000001400000027ffffffec00000014000000280;
		6'b001011:	xpb = 256'h000002c0000000000000016000000160000002bffffffea000000160000002c0;
		6'b001100:	xpb = 256'h00000300000000000000018000000180000002fffffffe800000018000000300;
		6'b001101:	xpb = 256'h0000034000000000000001a0000001a00000033ffffffe60000001a000000340;
		6'b001110:	xpb = 256'h0000038000000000000001c0000001c00000037ffffffe40000001c000000380;
		6'b001111:	xpb = 256'h000003c000000000000001e0000001e0000003bffffffe20000001e0000003c0;
		6'b010000:	xpb = 256'h00000400000000000000020000000200000003fffffffe000000020000000400;
		6'b010001:	xpb = 256'h000004400000000000000220000002200000043ffffffde00000022000000440;
		6'b010010:	xpb = 256'h000004800000000000000240000002400000047ffffffdc00000024000000480;
		6'b010011:	xpb = 256'h000004c0000000000000026000000260000004bffffffda000000260000004c0;
		6'b010100:	xpb = 256'h00000500000000000000028000000280000004fffffffd800000028000000500;
		6'b010101:	xpb = 256'h0000054000000000000002a0000002a00000053ffffffd60000002a000000540;
		6'b010110:	xpb = 256'h0000058000000000000002c0000002c00000057ffffffd40000002c000000580;
		6'b010111:	xpb = 256'h000005c000000000000002e0000002e0000005bffffffd20000002e0000005c0;
		6'b011000:	xpb = 256'h00000600000000000000030000000300000005fffffffd000000030000000600;
		6'b011001:	xpb = 256'h000006400000000000000320000003200000063ffffffce00000032000000640;
		6'b011010:	xpb = 256'h000006800000000000000340000003400000067ffffffcc00000034000000680;
		6'b011011:	xpb = 256'h000006c0000000000000036000000360000006bffffffca000000360000006c0;
		6'b011100:	xpb = 256'h00000700000000000000038000000380000006fffffffc800000038000000700;
		6'b011101:	xpb = 256'h0000074000000000000003a0000003a00000073ffffffc60000003a000000740;
		6'b011110:	xpb = 256'h0000078000000000000003c0000003c00000077ffffffc40000003c000000780;
		6'b011111:	xpb = 256'h000007c000000000000003e0000003e0000007bffffffc20000003e0000007c0;
		6'b100000:	xpb = 256'h00000800000000000000040000000400000007fffffffc000000040000000800;
		6'b100001:	xpb = 256'h000008400000000000000420000004200000083ffffffbe00000042000000840;
		6'b100010:	xpb = 256'h000008800000000000000440000004400000087ffffffbc00000044000000880;
		6'b100011:	xpb = 256'h000008c0000000000000046000000460000008bffffffba000000460000008c0;
		6'b100100:	xpb = 256'h00000900000000000000048000000480000008fffffffb800000048000000900;
		6'b100101:	xpb = 256'h0000094000000000000004a0000004a00000093ffffffb60000004a000000940;
		6'b100110:	xpb = 256'h0000098000000000000004c0000004c00000097ffffffb40000004c000000980;
		6'b100111:	xpb = 256'h000009c000000000000004e0000004e0000009bffffffb20000004e0000009c0;
		6'b101000:	xpb = 256'h00000a00000000000000050000000500000009fffffffb000000050000000a00;
		6'b101001:	xpb = 256'h00000a4000000000000005200000052000000a3ffffffae00000052000000a40;
		6'b101010:	xpb = 256'h00000a8000000000000005400000054000000a7ffffffac00000054000000a80;
		6'b101011:	xpb = 256'h00000ac000000000000005600000056000000abffffffaa00000056000000ac0;
		6'b101100:	xpb = 256'h00000b0000000000000005800000058000000afffffffa800000058000000b00;
		6'b101101:	xpb = 256'h00000b4000000000000005a0000005a000000b3ffffffa60000005a000000b40;
		6'b101110:	xpb = 256'h00000b8000000000000005c0000005c000000b7ffffffa40000005c000000b80;
		6'b101111:	xpb = 256'h00000bc000000000000005e0000005e000000bbffffffa20000005e000000bc0;
		6'b110000:	xpb = 256'h00000c0000000000000006000000060000000bfffffffa000000060000000c00;
		6'b110001:	xpb = 256'h00000c4000000000000006200000062000000c3ffffff9e00000062000000c40;
		6'b110010:	xpb = 256'h00000c8000000000000006400000064000000c7ffffff9c00000064000000c80;
		6'b110011:	xpb = 256'h00000cc000000000000006600000066000000cbffffff9a00000066000000cc0;
		6'b110100:	xpb = 256'h00000d0000000000000006800000068000000cfffffff9800000068000000d00;
		6'b110101:	xpb = 256'h00000d4000000000000006a0000006a000000d3ffffff960000006a000000d40;
		6'b110110:	xpb = 256'h00000d8000000000000006c0000006c000000d7ffffff940000006c000000d80;
		6'b110111:	xpb = 256'h00000dc000000000000006e0000006e000000dbffffff920000006e000000dc0;
		6'b111000:	xpb = 256'h00000e0000000000000007000000070000000dfffffff9000000070000000e00;
		6'b111001:	xpb = 256'h00000e4000000000000007200000072000000e3ffffff8e00000072000000e40;
		6'b111010:	xpb = 256'h00000e8000000000000007400000074000000e7ffffff8c00000074000000e80;
		6'b111011:	xpb = 256'h00000ec000000000000007600000076000000ebffffff8a00000076000000ec0;
		6'b111100:	xpb = 256'h00000f0000000000000007800000078000000efffffff8800000078000000f00;
		6'b111101:	xpb = 256'h00000f4000000000000007a0000007a000000f3ffffff860000007a000000f40;
		6'b111110:	xpb = 256'h00000f8000000000000007c0000007c000000f7ffffff840000007c000000f80;
		6'b111111:	xpb = 256'h00000fc000000000000007e0000007e000000fbffffff820000007e000000fc0;
	endcase
end
endmodule

module xpb_26_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000100000000000000008000000080000000ffffffff8000000080000001000;
		6'b000010:	xpb = 256'h0000200000000000000010000000100000001ffffffff0000000100000002000;
		6'b000011:	xpb = 256'h0000300000000000000018000000180000002fffffffe8000000180000003000;
		6'b000100:	xpb = 256'h0000400000000000000020000000200000003fffffffe0000000200000004000;
		6'b000101:	xpb = 256'h0000500000000000000028000000280000004fffffffd8000000280000005000;
		6'b000110:	xpb = 256'h0000600000000000000030000000300000005fffffffd0000000300000006000;
		6'b000111:	xpb = 256'h0000700000000000000038000000380000006fffffffc8000000380000007000;
		6'b001000:	xpb = 256'h0000800000000000000040000000400000007fffffffc0000000400000008000;
		6'b001001:	xpb = 256'h0000900000000000000048000000480000008fffffffb8000000480000009000;
		6'b001010:	xpb = 256'h0000a00000000000000050000000500000009fffffffb000000050000000a000;
		6'b001011:	xpb = 256'h0000b0000000000000005800000058000000afffffffa800000058000000b000;
		6'b001100:	xpb = 256'h0000c0000000000000006000000060000000bfffffffa000000060000000c000;
		6'b001101:	xpb = 256'h0000d0000000000000006800000068000000cfffffff9800000068000000d000;
		6'b001110:	xpb = 256'h0000e0000000000000007000000070000000dfffffff9000000070000000e000;
		6'b001111:	xpb = 256'h0000f0000000000000007800000078000000efffffff8800000078000000f000;
		6'b010000:	xpb = 256'h000100000000000000008000000080000000ffffffff80000000800000010000;
		6'b010001:	xpb = 256'h0001100000000000000088000000880000010fffffff78000000880000011000;
		6'b010010:	xpb = 256'h0001200000000000000090000000900000011fffffff70000000900000012000;
		6'b010011:	xpb = 256'h0001300000000000000098000000980000012fffffff68000000980000013000;
		6'b010100:	xpb = 256'h00014000000000000000a0000000a00000013fffffff60000000a00000014000;
		6'b010101:	xpb = 256'h00015000000000000000a8000000a80000014fffffff58000000a80000015000;
		6'b010110:	xpb = 256'h00016000000000000000b0000000b00000015fffffff50000000b00000016000;
		6'b010111:	xpb = 256'h00017000000000000000b8000000b80000016fffffff48000000b80000017000;
		6'b011000:	xpb = 256'h00018000000000000000c0000000c00000017fffffff40000000c00000018000;
		6'b011001:	xpb = 256'h00019000000000000000c8000000c80000018fffffff38000000c80000019000;
		6'b011010:	xpb = 256'h0001a000000000000000d0000000d00000019fffffff30000000d0000001a000;
		6'b011011:	xpb = 256'h0001b000000000000000d8000000d8000001afffffff28000000d8000001b000;
		6'b011100:	xpb = 256'h0001c000000000000000e0000000e0000001bfffffff20000000e0000001c000;
		6'b011101:	xpb = 256'h0001d000000000000000e8000000e8000001cfffffff18000000e8000001d000;
		6'b011110:	xpb = 256'h0001e000000000000000f0000000f0000001dfffffff10000000f0000001e000;
		6'b011111:	xpb = 256'h0001f000000000000000f8000000f8000001efffffff08000000f8000001f000;
		6'b100000:	xpb = 256'h000200000000000000010000000100000001ffffffff00000001000000020000;
		6'b100001:	xpb = 256'h0002100000000000000108000001080000020ffffffef8000001080000021000;
		6'b100010:	xpb = 256'h0002200000000000000110000001100000021ffffffef0000001100000022000;
		6'b100011:	xpb = 256'h0002300000000000000118000001180000022ffffffee8000001180000023000;
		6'b100100:	xpb = 256'h0002400000000000000120000001200000023ffffffee0000001200000024000;
		6'b100101:	xpb = 256'h0002500000000000000128000001280000024ffffffed8000001280000025000;
		6'b100110:	xpb = 256'h0002600000000000000130000001300000025ffffffed0000001300000026000;
		6'b100111:	xpb = 256'h0002700000000000000138000001380000026ffffffec8000001380000027000;
		6'b101000:	xpb = 256'h0002800000000000000140000001400000027ffffffec0000001400000028000;
		6'b101001:	xpb = 256'h0002900000000000000148000001480000028ffffffeb8000001480000029000;
		6'b101010:	xpb = 256'h0002a00000000000000150000001500000029ffffffeb000000150000002a000;
		6'b101011:	xpb = 256'h0002b0000000000000015800000158000002affffffea800000158000002b000;
		6'b101100:	xpb = 256'h0002c0000000000000016000000160000002bffffffea000000160000002c000;
		6'b101101:	xpb = 256'h0002d0000000000000016800000168000002cffffffe9800000168000002d000;
		6'b101110:	xpb = 256'h0002e0000000000000017000000170000002dffffffe9000000170000002e000;
		6'b101111:	xpb = 256'h0002f0000000000000017800000178000002effffffe8800000178000002f000;
		6'b110000:	xpb = 256'h000300000000000000018000000180000002fffffffe80000001800000030000;
		6'b110001:	xpb = 256'h0003100000000000000188000001880000030ffffffe78000001880000031000;
		6'b110010:	xpb = 256'h0003200000000000000190000001900000031ffffffe70000001900000032000;
		6'b110011:	xpb = 256'h0003300000000000000198000001980000032ffffffe68000001980000033000;
		6'b110100:	xpb = 256'h00034000000000000001a0000001a00000033ffffffe60000001a00000034000;
		6'b110101:	xpb = 256'h00035000000000000001a8000001a80000034ffffffe58000001a80000035000;
		6'b110110:	xpb = 256'h00036000000000000001b0000001b00000035ffffffe50000001b00000036000;
		6'b110111:	xpb = 256'h00037000000000000001b8000001b80000036ffffffe48000001b80000037000;
		6'b111000:	xpb = 256'h00038000000000000001c0000001c00000037ffffffe40000001c00000038000;
		6'b111001:	xpb = 256'h00039000000000000001c8000001c80000038ffffffe38000001c80000039000;
		6'b111010:	xpb = 256'h0003a000000000000001d0000001d00000039ffffffe30000001d0000003a000;
		6'b111011:	xpb = 256'h0003b000000000000001d8000001d8000003affffffe28000001d8000003b000;
		6'b111100:	xpb = 256'h0003c000000000000001e0000001e0000003bffffffe20000001e0000003c000;
		6'b111101:	xpb = 256'h0003d000000000000001e8000001e8000003cffffffe18000001e8000003d000;
		6'b111110:	xpb = 256'h0003e000000000000001f0000001f0000003dffffffe10000001f0000003e000;
		6'b111111:	xpb = 256'h0003f000000000000001f8000001f8000003effffffe08000001f8000003f000;
	endcase
end
endmodule

module xpb_27_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h000200000000000000010000000100000001ffffffff00000001000000020000;
		5'b00010:	xpb = 256'h000400000000000000020000000200000003fffffffe00000002000000040000;
		5'b00011:	xpb = 256'h000600000000000000030000000300000005fffffffd00000003000000060000;
		5'b00100:	xpb = 256'h000800000000000000040000000400000007fffffffc00000004000000080000;
		5'b00101:	xpb = 256'h000a00000000000000050000000500000009fffffffb000000050000000a0000;
		5'b00110:	xpb = 256'h000c0000000000000006000000060000000bfffffffa000000060000000c0000;
		5'b00111:	xpb = 256'h000e0000000000000007000000070000000dfffffff9000000070000000e0000;
		5'b01000:	xpb = 256'h00100000000000000008000000080000000ffffffff800000008000000100000;
		5'b01001:	xpb = 256'h001200000000000000090000000900000011fffffff700000009000000120000;
		5'b01010:	xpb = 256'h0014000000000000000a0000000a00000013fffffff60000000a000000140000;
		5'b01011:	xpb = 256'h0016000000000000000b0000000b00000015fffffff50000000b000000160000;
		5'b01100:	xpb = 256'h0018000000000000000c0000000c00000017fffffff40000000c000000180000;
		5'b01101:	xpb = 256'h001a000000000000000d0000000d00000019fffffff30000000d0000001a0000;
		5'b01110:	xpb = 256'h001c000000000000000e0000000e0000001bfffffff20000000e0000001c0000;
		5'b01111:	xpb = 256'h001e000000000000000f0000000f0000001dfffffff10000000f0000001e0000;
		5'b10000:	xpb = 256'h00200000000000000010000000100000001ffffffff000000010000000200000;
		5'b10001:	xpb = 256'h002200000000000000110000001100000021ffffffef00000011000000220000;
		5'b10010:	xpb = 256'h002400000000000000120000001200000023ffffffee00000012000000240000;
		5'b10011:	xpb = 256'h002600000000000000130000001300000025ffffffed00000013000000260000;
		5'b10100:	xpb = 256'h002800000000000000140000001400000027ffffffec00000014000000280000;
		5'b10101:	xpb = 256'h002a00000000000000150000001500000029ffffffeb000000150000002a0000;
		5'b10110:	xpb = 256'h002c0000000000000016000000160000002bffffffea000000160000002c0000;
		5'b10111:	xpb = 256'h002e0000000000000017000000170000002dffffffe9000000170000002e0000;
		5'b11000:	xpb = 256'h00300000000000000018000000180000002fffffffe800000018000000300000;
		5'b11001:	xpb = 256'h003200000000000000190000001900000031ffffffe700000019000000320000;
		5'b11010:	xpb = 256'h0034000000000000001a0000001a00000033ffffffe60000001a000000340000;
		5'b11011:	xpb = 256'h0036000000000000001b0000001b00000035ffffffe50000001b000000360000;
		5'b11100:	xpb = 256'h0038000000000000001c0000001c00000037ffffffe40000001c000000380000;
		5'b11101:	xpb = 256'h003a000000000000001d0000001d00000039ffffffe30000001d0000003a0000;
		5'b11110:	xpb = 256'h003c000000000000001e0000001e0000003bffffffe20000001e0000003c0000;
		5'b11111:	xpb = 256'h003e000000000000001f0000001f0000003dffffffe10000001f0000003e0000;
	endcase
end
endmodule

module xpb_27_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00400000000000000020000000200000003fffffffe000000020000000400000;
		6'b000010:	xpb = 256'h00800000000000000040000000400000007fffffffc000000040000000800000;
		6'b000011:	xpb = 256'h00c0000000000000006000000060000000bfffffffa000000060000000c00000;
		6'b000100:	xpb = 256'h0100000000000000008000000080000000ffffffff8000000080000001000000;
		6'b000101:	xpb = 256'h014000000000000000a0000000a00000013fffffff60000000a0000001400000;
		6'b000110:	xpb = 256'h018000000000000000c0000000c00000017fffffff40000000c0000001800000;
		6'b000111:	xpb = 256'h01c000000000000000e0000000e0000001bfffffff20000000e0000001c00000;
		6'b001000:	xpb = 256'h0200000000000000010000000100000001ffffffff0000000100000002000000;
		6'b001001:	xpb = 256'h02400000000000000120000001200000023ffffffee000000120000002400000;
		6'b001010:	xpb = 256'h02800000000000000140000001400000027ffffffec000000140000002800000;
		6'b001011:	xpb = 256'h02c0000000000000016000000160000002bffffffea000000160000002c00000;
		6'b001100:	xpb = 256'h0300000000000000018000000180000002fffffffe8000000180000003000000;
		6'b001101:	xpb = 256'h034000000000000001a0000001a00000033ffffffe60000001a0000003400000;
		6'b001110:	xpb = 256'h038000000000000001c0000001c00000037ffffffe40000001c0000003800000;
		6'b001111:	xpb = 256'h03c000000000000001e0000001e0000003bffffffe20000001e0000003c00000;
		6'b010000:	xpb = 256'h0400000000000000020000000200000003fffffffe0000000200000004000000;
		6'b010001:	xpb = 256'h04400000000000000220000002200000043ffffffde000000220000004400000;
		6'b010010:	xpb = 256'h04800000000000000240000002400000047ffffffdc000000240000004800000;
		6'b010011:	xpb = 256'h04c0000000000000026000000260000004bffffffda000000260000004c00000;
		6'b010100:	xpb = 256'h0500000000000000028000000280000004fffffffd8000000280000005000000;
		6'b010101:	xpb = 256'h054000000000000002a0000002a00000053ffffffd60000002a0000005400000;
		6'b010110:	xpb = 256'h058000000000000002c0000002c00000057ffffffd40000002c0000005800000;
		6'b010111:	xpb = 256'h05c000000000000002e0000002e0000005bffffffd20000002e0000005c00000;
		6'b011000:	xpb = 256'h0600000000000000030000000300000005fffffffd0000000300000006000000;
		6'b011001:	xpb = 256'h06400000000000000320000003200000063ffffffce000000320000006400000;
		6'b011010:	xpb = 256'h06800000000000000340000003400000067ffffffcc000000340000006800000;
		6'b011011:	xpb = 256'h06c0000000000000036000000360000006bffffffca000000360000006c00000;
		6'b011100:	xpb = 256'h0700000000000000038000000380000006fffffffc8000000380000007000000;
		6'b011101:	xpb = 256'h074000000000000003a0000003a00000073ffffffc60000003a0000007400000;
		6'b011110:	xpb = 256'h078000000000000003c0000003c00000077ffffffc40000003c0000007800000;
		6'b011111:	xpb = 256'h07c000000000000003e0000003e0000007bffffffc20000003e0000007c00000;
		6'b100000:	xpb = 256'h0800000000000000040000000400000007fffffffc0000000400000008000000;
		6'b100001:	xpb = 256'h08400000000000000420000004200000083ffffffbe000000420000008400000;
		6'b100010:	xpb = 256'h08800000000000000440000004400000087ffffffbc000000440000008800000;
		6'b100011:	xpb = 256'h08c0000000000000046000000460000008bffffffba000000460000008c00000;
		6'b100100:	xpb = 256'h0900000000000000048000000480000008fffffffb8000000480000009000000;
		6'b100101:	xpb = 256'h094000000000000004a0000004a00000093ffffffb60000004a0000009400000;
		6'b100110:	xpb = 256'h098000000000000004c0000004c00000097ffffffb40000004c0000009800000;
		6'b100111:	xpb = 256'h09c000000000000004e0000004e0000009bffffffb20000004e0000009c00000;
		6'b101000:	xpb = 256'h0a00000000000000050000000500000009fffffffb000000050000000a000000;
		6'b101001:	xpb = 256'h0a4000000000000005200000052000000a3ffffffae00000052000000a400000;
		6'b101010:	xpb = 256'h0a8000000000000005400000054000000a7ffffffac00000054000000a800000;
		6'b101011:	xpb = 256'h0ac000000000000005600000056000000abffffffaa00000056000000ac00000;
		6'b101100:	xpb = 256'h0b0000000000000005800000058000000afffffffa800000058000000b000000;
		6'b101101:	xpb = 256'h0b4000000000000005a0000005a000000b3ffffffa60000005a000000b400000;
		6'b101110:	xpb = 256'h0b8000000000000005c0000005c000000b7ffffffa40000005c000000b800000;
		6'b101111:	xpb = 256'h0bc000000000000005e0000005e000000bbffffffa20000005e000000bc00000;
		6'b110000:	xpb = 256'h0c0000000000000006000000060000000bfffffffa000000060000000c000000;
		6'b110001:	xpb = 256'h0c4000000000000006200000062000000c3ffffff9e00000062000000c400000;
		6'b110010:	xpb = 256'h0c8000000000000006400000064000000c7ffffff9c00000064000000c800000;
		6'b110011:	xpb = 256'h0cc000000000000006600000066000000cbffffff9a00000066000000cc00000;
		6'b110100:	xpb = 256'h0d0000000000000006800000068000000cfffffff9800000068000000d000000;
		6'b110101:	xpb = 256'h0d4000000000000006a0000006a000000d3ffffff960000006a000000d400000;
		6'b110110:	xpb = 256'h0d8000000000000006c0000006c000000d7ffffff940000006c000000d800000;
		6'b110111:	xpb = 256'h0dc000000000000006e0000006e000000dbffffff920000006e000000dc00000;
		6'b111000:	xpb = 256'h0e0000000000000007000000070000000dfffffff9000000070000000e000000;
		6'b111001:	xpb = 256'h0e4000000000000007200000072000000e3ffffff8e00000072000000e400000;
		6'b111010:	xpb = 256'h0e8000000000000007400000074000000e7ffffff8c00000074000000e800000;
		6'b111011:	xpb = 256'h0ec000000000000007600000076000000ebffffff8a00000076000000ec00000;
		6'b111100:	xpb = 256'h0f0000000000000007800000078000000efffffff8800000078000000f000000;
		6'b111101:	xpb = 256'h0f4000000000000007a0000007a000000f3ffffff860000007a000000f400000;
		6'b111110:	xpb = 256'h0f8000000000000007c0000007c000000f7ffffff840000007c000000f800000;
		6'b111111:	xpb = 256'h0fc000000000000007e0000007e000000fbffffff820000007e000000fc00000;
	endcase
end
endmodule

module xpb_27_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h100000000000000008000000080000000ffffffff80000000800000010000000;
		6'b000010:	xpb = 256'h200000000000000010000000100000001ffffffff00000001000000020000000;
		6'b000011:	xpb = 256'h300000000000000018000000180000002fffffffe80000001800000030000000;
		6'b000100:	xpb = 256'h400000000000000020000000200000003fffffffe00000002000000040000000;
		6'b000101:	xpb = 256'h500000000000000028000000280000004fffffffd80000002800000050000000;
		6'b000110:	xpb = 256'h600000000000000030000000300000005fffffffd00000003000000060000000;
		6'b000111:	xpb = 256'h700000000000000038000000380000006fffffffc80000003800000070000000;
		6'b001000:	xpb = 256'h800000000000000040000000400000007fffffffc00000004000000080000000;
		6'b001001:	xpb = 256'h900000000000000048000000480000008fffffffb80000004800000090000000;
		6'b001010:	xpb = 256'ha00000000000000050000000500000009fffffffb000000050000000a0000000;
		6'b001011:	xpb = 256'hb0000000000000005800000058000000afffffffa800000058000000b0000000;
		6'b001100:	xpb = 256'hc0000000000000006000000060000000bfffffffa000000060000000c0000000;
		6'b001101:	xpb = 256'hd0000000000000006800000068000000cfffffff9800000068000000d0000000;
		6'b001110:	xpb = 256'he0000000000000007000000070000000dfffffff9000000070000000e0000000;
		6'b001111:	xpb = 256'hf0000000000000007800000078000000efffffff8800000078000000f0000000;
		6'b010000:	xpb = 256'h00000001000000008000000080000001000000007fffffff8000000100000001;
		6'b010001:	xpb = 256'h100000010000000088000000880000011000000077ffffff8800000110000001;
		6'b010010:	xpb = 256'h20000001000000009000000090000001200000006fffffff9000000120000001;
		6'b010011:	xpb = 256'h300000010000000098000000980000013000000067ffffff9800000130000001;
		6'b010100:	xpb = 256'h4000000100000000a0000000a0000001400000005fffffffa000000140000001;
		6'b010101:	xpb = 256'h5000000100000000a8000000a80000015000000057ffffffa800000150000001;
		6'b010110:	xpb = 256'h6000000100000000b0000000b0000001600000004fffffffb000000160000001;
		6'b010111:	xpb = 256'h7000000100000000b8000000b80000017000000047ffffffb800000170000001;
		6'b011000:	xpb = 256'h8000000100000000c0000000c0000001800000003fffffffc000000180000001;
		6'b011001:	xpb = 256'h9000000100000000c8000000c80000019000000037ffffffc800000190000001;
		6'b011010:	xpb = 256'ha000000100000000d0000000d0000001a00000002fffffffd0000001a0000001;
		6'b011011:	xpb = 256'hb000000100000000d8000000d8000001b000000027ffffffd8000001b0000001;
		6'b011100:	xpb = 256'hc000000100000000e0000000e0000001c00000001fffffffe0000001c0000001;
		6'b011101:	xpb = 256'hd000000100000000e8000000e8000001d000000017ffffffe8000001d0000001;
		6'b011110:	xpb = 256'he000000100000000f0000000f0000001e00000000ffffffff0000001e0000001;
		6'b011111:	xpb = 256'hf000000100000000f8000000f8000001f000000007fffffff8000001f0000001;
		6'b100000:	xpb = 256'h0000000200000001000000010000000200000000ffffffff0000000200000002;
		6'b100001:	xpb = 256'h1000000200000001080000010800000210000000f7ffffff0800000210000002;
		6'b100010:	xpb = 256'h2000000200000001100000011000000220000000efffffff1000000220000002;
		6'b100011:	xpb = 256'h3000000200000001180000011800000230000000e7ffffff1800000230000002;
		6'b100100:	xpb = 256'h4000000200000001200000012000000240000000dfffffff2000000240000002;
		6'b100101:	xpb = 256'h5000000200000001280000012800000250000000d7ffffff2800000250000002;
		6'b100110:	xpb = 256'h6000000200000001300000013000000260000000cfffffff3000000260000002;
		6'b100111:	xpb = 256'h7000000200000001380000013800000270000000c7ffffff3800000270000002;
		6'b101000:	xpb = 256'h8000000200000001400000014000000280000000bfffffff4000000280000002;
		6'b101001:	xpb = 256'h9000000200000001480000014800000290000000b7ffffff4800000290000002;
		6'b101010:	xpb = 256'ha0000002000000015000000150000002a0000000afffffff50000002a0000002;
		6'b101011:	xpb = 256'hb0000002000000015800000158000002b0000000a7ffffff58000002b0000002;
		6'b101100:	xpb = 256'hc0000002000000016000000160000002c00000009fffffff60000002c0000002;
		6'b101101:	xpb = 256'hd0000002000000016800000168000002d000000097ffffff68000002d0000002;
		6'b101110:	xpb = 256'he0000002000000017000000170000002e00000008fffffff70000002e0000002;
		6'b101111:	xpb = 256'hf0000002000000017800000178000002f000000087ffffff78000002f0000002;
		6'b110000:	xpb = 256'h00000003000000018000000180000003000000017ffffffe8000000300000003;
		6'b110001:	xpb = 256'h100000030000000188000001880000031000000177fffffe8800000310000003;
		6'b110010:	xpb = 256'h20000003000000019000000190000003200000016ffffffe9000000320000003;
		6'b110011:	xpb = 256'h300000030000000198000001980000033000000167fffffe9800000330000003;
		6'b110100:	xpb = 256'h4000000300000001a0000001a0000003400000015ffffffea000000340000003;
		6'b110101:	xpb = 256'h5000000300000001a8000001a80000035000000157fffffea800000350000003;
		6'b110110:	xpb = 256'h6000000300000001b0000001b0000003600000014ffffffeb000000360000003;
		6'b110111:	xpb = 256'h7000000300000001b8000001b80000037000000147fffffeb800000370000003;
		6'b111000:	xpb = 256'h8000000300000001c0000001c0000003800000013ffffffec000000380000003;
		6'b111001:	xpb = 256'h9000000300000001c8000001c80000039000000137fffffec800000390000003;
		6'b111010:	xpb = 256'ha000000300000001d0000001d0000003a00000012ffffffed0000003a0000003;
		6'b111011:	xpb = 256'hb000000300000001d8000001d8000003b000000127fffffed8000003b0000003;
		6'b111100:	xpb = 256'hc000000300000001e0000001e0000003c00000011ffffffee0000003c0000003;
		6'b111101:	xpb = 256'hd000000300000001e8000001e8000003d000000117fffffee8000003d0000003;
		6'b111110:	xpb = 256'he000000300000001f0000001f0000003e00000010ffffffef0000003e0000003;
		6'b111111:	xpb = 256'hf000000300000001f8000001f8000003f000000107fffffef8000003f0000003;
	endcase
end
endmodule

module xpb_28_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000200000001000000010000000200000000ffffffff0000000200000002;
		5'b00010:	xpb = 256'h0000000400000002000000020000000400000001fffffffe0000000400000004;
		5'b00011:	xpb = 256'h0000000600000003000000030000000600000002fffffffd0000000600000006;
		5'b00100:	xpb = 256'h0000000800000004000000040000000800000003fffffffc0000000800000008;
		5'b00101:	xpb = 256'h0000000a00000005000000050000000a00000004fffffffb0000000a0000000a;
		5'b00110:	xpb = 256'h0000000c00000006000000060000000c00000005fffffffa0000000c0000000c;
		5'b00111:	xpb = 256'h0000000e00000007000000070000000e00000006fffffff90000000e0000000e;
		5'b01000:	xpb = 256'h0000001000000008000000080000001000000007fffffff80000001000000010;
		5'b01001:	xpb = 256'h0000001200000009000000090000001200000008fffffff70000001200000012;
		5'b01010:	xpb = 256'h000000140000000a0000000a0000001400000009fffffff60000001400000014;
		5'b01011:	xpb = 256'h000000160000000b0000000b000000160000000afffffff50000001600000016;
		5'b01100:	xpb = 256'h000000180000000c0000000c000000180000000bfffffff40000001800000018;
		5'b01101:	xpb = 256'h0000001a0000000d0000000d0000001a0000000cfffffff30000001a0000001a;
		5'b01110:	xpb = 256'h0000001c0000000e0000000e0000001c0000000dfffffff20000001c0000001c;
		5'b01111:	xpb = 256'h0000001e0000000f0000000f0000001e0000000efffffff10000001e0000001e;
		5'b10000:	xpb = 256'h000000200000001000000010000000200000000ffffffff00000002000000020;
		5'b10001:	xpb = 256'h0000002200000011000000110000002200000010ffffffef0000002200000022;
		5'b10010:	xpb = 256'h0000002400000012000000120000002400000011ffffffee0000002400000024;
		5'b10011:	xpb = 256'h0000002600000013000000130000002600000012ffffffed0000002600000026;
		5'b10100:	xpb = 256'h0000002800000014000000140000002800000013ffffffec0000002800000028;
		5'b10101:	xpb = 256'h0000002a00000015000000150000002a00000014ffffffeb0000002a0000002a;
		5'b10110:	xpb = 256'h0000002c00000016000000160000002c00000015ffffffea0000002c0000002c;
		5'b10111:	xpb = 256'h0000002e00000017000000170000002e00000016ffffffe90000002e0000002e;
		5'b11000:	xpb = 256'h0000003000000018000000180000003000000017ffffffe80000003000000030;
		5'b11001:	xpb = 256'h0000003200000019000000190000003200000018ffffffe70000003200000032;
		5'b11010:	xpb = 256'h000000340000001a0000001a0000003400000019ffffffe60000003400000034;
		5'b11011:	xpb = 256'h000000360000001b0000001b000000360000001affffffe50000003600000036;
		5'b11100:	xpb = 256'h000000380000001c0000001c000000380000001bffffffe40000003800000038;
		5'b11101:	xpb = 256'h0000003a0000001d0000001d0000003a0000001cffffffe30000003a0000003a;
		5'b11110:	xpb = 256'h0000003c0000001e0000001e0000003c0000001dffffffe20000003c0000003c;
		5'b11111:	xpb = 256'h0000003e0000001f0000001f0000003e0000001effffffe10000003e0000003e;
	endcase
end
endmodule

module xpb_28_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h000000400000002000000020000000400000001fffffffe00000004000000040;
		6'b000010:	xpb = 256'h000000800000004000000040000000800000003fffffffc00000008000000080;
		6'b000011:	xpb = 256'h000000c00000006000000060000000c00000005fffffffa0000000c0000000c0;
		6'b000100:	xpb = 256'h000001000000008000000080000001000000007fffffff800000010000000100;
		6'b000101:	xpb = 256'h00000140000000a0000000a0000001400000009fffffff600000014000000140;
		6'b000110:	xpb = 256'h00000180000000c0000000c000000180000000bfffffff400000018000000180;
		6'b000111:	xpb = 256'h000001c0000000e0000000e0000001c0000000dfffffff20000001c0000001c0;
		6'b001000:	xpb = 256'h00000200000001000000010000000200000000ffffffff000000020000000200;
		6'b001001:	xpb = 256'h000002400000012000000120000002400000011ffffffee00000024000000240;
		6'b001010:	xpb = 256'h000002800000014000000140000002800000013ffffffec00000028000000280;
		6'b001011:	xpb = 256'h000002c00000016000000160000002c00000015ffffffea0000002c0000002c0;
		6'b001100:	xpb = 256'h000003000000018000000180000003000000017ffffffe800000030000000300;
		6'b001101:	xpb = 256'h00000340000001a0000001a0000003400000019ffffffe600000034000000340;
		6'b001110:	xpb = 256'h00000380000001c0000001c000000380000001bffffffe400000038000000380;
		6'b001111:	xpb = 256'h000003c0000001e0000001e0000003c0000001dffffffe20000003c0000003c0;
		6'b010000:	xpb = 256'h00000400000002000000020000000400000001fffffffe000000040000000400;
		6'b010001:	xpb = 256'h000004400000022000000220000004400000021ffffffde00000044000000440;
		6'b010010:	xpb = 256'h000004800000024000000240000004800000023ffffffdc00000048000000480;
		6'b010011:	xpb = 256'h000004c00000026000000260000004c00000025ffffffda0000004c0000004c0;
		6'b010100:	xpb = 256'h000005000000028000000280000005000000027ffffffd800000050000000500;
		6'b010101:	xpb = 256'h00000540000002a0000002a0000005400000029ffffffd600000054000000540;
		6'b010110:	xpb = 256'h00000580000002c0000002c000000580000002bffffffd400000058000000580;
		6'b010111:	xpb = 256'h000005c0000002e0000002e0000005c0000002dffffffd20000005c0000005c0;
		6'b011000:	xpb = 256'h00000600000003000000030000000600000002fffffffd000000060000000600;
		6'b011001:	xpb = 256'h000006400000032000000320000006400000031ffffffce00000064000000640;
		6'b011010:	xpb = 256'h000006800000034000000340000006800000033ffffffcc00000068000000680;
		6'b011011:	xpb = 256'h000006c00000036000000360000006c00000035ffffffca0000006c0000006c0;
		6'b011100:	xpb = 256'h000007000000038000000380000007000000037ffffffc800000070000000700;
		6'b011101:	xpb = 256'h00000740000003a0000003a0000007400000039ffffffc600000074000000740;
		6'b011110:	xpb = 256'h00000780000003c0000003c000000780000003bffffffc400000078000000780;
		6'b011111:	xpb = 256'h000007c0000003e0000003e0000007c0000003dffffffc20000007c0000007c0;
		6'b100000:	xpb = 256'h00000800000004000000040000000800000003fffffffc000000080000000800;
		6'b100001:	xpb = 256'h000008400000042000000420000008400000041ffffffbe00000084000000840;
		6'b100010:	xpb = 256'h000008800000044000000440000008800000043ffffffbc00000088000000880;
		6'b100011:	xpb = 256'h000008c00000046000000460000008c00000045ffffffba0000008c0000008c0;
		6'b100100:	xpb = 256'h000009000000048000000480000009000000047ffffffb800000090000000900;
		6'b100101:	xpb = 256'h00000940000004a0000004a0000009400000049ffffffb600000094000000940;
		6'b100110:	xpb = 256'h00000980000004c0000004c000000980000004bffffffb400000098000000980;
		6'b100111:	xpb = 256'h000009c0000004e0000004e0000009c0000004dffffffb20000009c0000009c0;
		6'b101000:	xpb = 256'h00000a00000005000000050000000a00000004fffffffb0000000a0000000a00;
		6'b101001:	xpb = 256'h00000a40000005200000052000000a400000051ffffffae000000a4000000a40;
		6'b101010:	xpb = 256'h00000a80000005400000054000000a800000053ffffffac000000a8000000a80;
		6'b101011:	xpb = 256'h00000ac0000005600000056000000ac00000055ffffffaa000000ac000000ac0;
		6'b101100:	xpb = 256'h00000b00000005800000058000000b000000057ffffffa8000000b0000000b00;
		6'b101101:	xpb = 256'h00000b40000005a0000005a000000b400000059ffffffa6000000b4000000b40;
		6'b101110:	xpb = 256'h00000b80000005c0000005c000000b80000005bffffffa4000000b8000000b80;
		6'b101111:	xpb = 256'h00000bc0000005e0000005e000000bc0000005dffffffa2000000bc000000bc0;
		6'b110000:	xpb = 256'h00000c00000006000000060000000c00000005fffffffa0000000c0000000c00;
		6'b110001:	xpb = 256'h00000c40000006200000062000000c400000061ffffff9e000000c4000000c40;
		6'b110010:	xpb = 256'h00000c80000006400000064000000c800000063ffffff9c000000c8000000c80;
		6'b110011:	xpb = 256'h00000cc0000006600000066000000cc00000065ffffff9a000000cc000000cc0;
		6'b110100:	xpb = 256'h00000d00000006800000068000000d000000067ffffff98000000d0000000d00;
		6'b110101:	xpb = 256'h00000d40000006a0000006a000000d400000069ffffff96000000d4000000d40;
		6'b110110:	xpb = 256'h00000d80000006c0000006c000000d80000006bffffff94000000d8000000d80;
		6'b110111:	xpb = 256'h00000dc0000006e0000006e000000dc0000006dffffff92000000dc000000dc0;
		6'b111000:	xpb = 256'h00000e00000007000000070000000e00000006fffffff90000000e0000000e00;
		6'b111001:	xpb = 256'h00000e40000007200000072000000e400000071ffffff8e000000e4000000e40;
		6'b111010:	xpb = 256'h00000e80000007400000074000000e800000073ffffff8c000000e8000000e80;
		6'b111011:	xpb = 256'h00000ec0000007600000076000000ec00000075ffffff8a000000ec000000ec0;
		6'b111100:	xpb = 256'h00000f00000007800000078000000f000000077ffffff88000000f0000000f00;
		6'b111101:	xpb = 256'h00000f40000007a0000007a000000f400000079ffffff86000000f4000000f40;
		6'b111110:	xpb = 256'h00000f80000007c0000007c000000f80000007bffffff84000000f8000000f80;
		6'b111111:	xpb = 256'h00000fc0000007e0000007e000000fc0000007dffffff82000000fc000000fc0;
	endcase
end
endmodule

module xpb_28_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00001000000008000000080000001000000007fffffff8000000100000001000;
		6'b000010:	xpb = 256'h0000200000001000000010000000200000000ffffffff0000000200000002000;
		6'b000011:	xpb = 256'h00003000000018000000180000003000000017ffffffe8000000300000003000;
		6'b000100:	xpb = 256'h0000400000002000000020000000400000001fffffffe0000000400000004000;
		6'b000101:	xpb = 256'h00005000000028000000280000005000000027ffffffd8000000500000005000;
		6'b000110:	xpb = 256'h0000600000003000000030000000600000002fffffffd0000000600000006000;
		6'b000111:	xpb = 256'h00007000000038000000380000007000000037ffffffc8000000700000007000;
		6'b001000:	xpb = 256'h0000800000004000000040000000800000003fffffffc0000000800000008000;
		6'b001001:	xpb = 256'h00009000000048000000480000009000000047ffffffb8000000900000009000;
		6'b001010:	xpb = 256'h0000a00000005000000050000000a00000004fffffffb0000000a0000000a000;
		6'b001011:	xpb = 256'h0000b00000005800000058000000b000000057ffffffa8000000b0000000b000;
		6'b001100:	xpb = 256'h0000c00000006000000060000000c00000005fffffffa0000000c0000000c000;
		6'b001101:	xpb = 256'h0000d00000006800000068000000d000000067ffffff98000000d0000000d000;
		6'b001110:	xpb = 256'h0000e00000007000000070000000e00000006fffffff90000000e0000000e000;
		6'b001111:	xpb = 256'h0000f00000007800000078000000f000000077ffffff88000000f0000000f000;
		6'b010000:	xpb = 256'h0001000000008000000080000001000000007fffffff80000001000000010000;
		6'b010001:	xpb = 256'h00011000000088000000880000011000000087ffffff78000001100000011000;
		6'b010010:	xpb = 256'h0001200000009000000090000001200000008fffffff70000001200000012000;
		6'b010011:	xpb = 256'h00013000000098000000980000013000000097ffffff68000001300000013000;
		6'b010100:	xpb = 256'h000140000000a0000000a0000001400000009fffffff60000001400000014000;
		6'b010101:	xpb = 256'h000150000000a8000000a800000150000000a7ffffff58000001500000015000;
		6'b010110:	xpb = 256'h000160000000b0000000b000000160000000afffffff50000001600000016000;
		6'b010111:	xpb = 256'h000170000000b8000000b800000170000000b7ffffff48000001700000017000;
		6'b011000:	xpb = 256'h000180000000c0000000c000000180000000bfffffff40000001800000018000;
		6'b011001:	xpb = 256'h000190000000c8000000c800000190000000c7ffffff38000001900000019000;
		6'b011010:	xpb = 256'h0001a0000000d0000000d0000001a0000000cfffffff30000001a0000001a000;
		6'b011011:	xpb = 256'h0001b0000000d8000000d8000001b0000000d7ffffff28000001b0000001b000;
		6'b011100:	xpb = 256'h0001c0000000e0000000e0000001c0000000dfffffff20000001c0000001c000;
		6'b011101:	xpb = 256'h0001d0000000e8000000e8000001d0000000e7ffffff18000001d0000001d000;
		6'b011110:	xpb = 256'h0001e0000000f0000000f0000001e0000000efffffff10000001e0000001e000;
		6'b011111:	xpb = 256'h0001f0000000f8000000f8000001f0000000f7ffffff08000001f0000001f000;
		6'b100000:	xpb = 256'h000200000001000000010000000200000000ffffffff00000002000000020000;
		6'b100001:	xpb = 256'h00021000000108000001080000021000000107fffffef8000002100000021000;
		6'b100010:	xpb = 256'h0002200000011000000110000002200000010ffffffef0000002200000022000;
		6'b100011:	xpb = 256'h00023000000118000001180000023000000117fffffee8000002300000023000;
		6'b100100:	xpb = 256'h0002400000012000000120000002400000011ffffffee0000002400000024000;
		6'b100101:	xpb = 256'h00025000000128000001280000025000000127fffffed8000002500000025000;
		6'b100110:	xpb = 256'h0002600000013000000130000002600000012ffffffed0000002600000026000;
		6'b100111:	xpb = 256'h00027000000138000001380000027000000137fffffec8000002700000027000;
		6'b101000:	xpb = 256'h0002800000014000000140000002800000013ffffffec0000002800000028000;
		6'b101001:	xpb = 256'h00029000000148000001480000029000000147fffffeb8000002900000029000;
		6'b101010:	xpb = 256'h0002a00000015000000150000002a00000014ffffffeb0000002a0000002a000;
		6'b101011:	xpb = 256'h0002b00000015800000158000002b000000157fffffea8000002b0000002b000;
		6'b101100:	xpb = 256'h0002c00000016000000160000002c00000015ffffffea0000002c0000002c000;
		6'b101101:	xpb = 256'h0002d00000016800000168000002d000000167fffffe98000002d0000002d000;
		6'b101110:	xpb = 256'h0002e00000017000000170000002e00000016ffffffe90000002e0000002e000;
		6'b101111:	xpb = 256'h0002f00000017800000178000002f000000177fffffe88000002f0000002f000;
		6'b110000:	xpb = 256'h0003000000018000000180000003000000017ffffffe80000003000000030000;
		6'b110001:	xpb = 256'h00031000000188000001880000031000000187fffffe78000003100000031000;
		6'b110010:	xpb = 256'h0003200000019000000190000003200000018ffffffe70000003200000032000;
		6'b110011:	xpb = 256'h00033000000198000001980000033000000197fffffe68000003300000033000;
		6'b110100:	xpb = 256'h000340000001a0000001a0000003400000019ffffffe60000003400000034000;
		6'b110101:	xpb = 256'h000350000001a8000001a800000350000001a7fffffe58000003500000035000;
		6'b110110:	xpb = 256'h000360000001b0000001b000000360000001affffffe50000003600000036000;
		6'b110111:	xpb = 256'h000370000001b8000001b800000370000001b7fffffe48000003700000037000;
		6'b111000:	xpb = 256'h000380000001c0000001c000000380000001bffffffe40000003800000038000;
		6'b111001:	xpb = 256'h000390000001c8000001c800000390000001c7fffffe38000003900000039000;
		6'b111010:	xpb = 256'h0003a0000001d0000001d0000003a0000001cffffffe30000003a0000003a000;
		6'b111011:	xpb = 256'h0003b0000001d8000001d8000003b0000001d7fffffe28000003b0000003b000;
		6'b111100:	xpb = 256'h0003c0000001e0000001e0000003c0000001dffffffe20000003c0000003c000;
		6'b111101:	xpb = 256'h0003d0000001e8000001e8000003d0000001e7fffffe18000003d0000003d000;
		6'b111110:	xpb = 256'h0003e0000001f0000001f0000003e0000001effffffe10000003e0000003e000;
		6'b111111:	xpb = 256'h0003f0000001f8000001f8000003f0000001f7fffffe08000003f0000003f000;
	endcase
end
endmodule

module xpb_29_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h000200000001000000010000000200000000ffffffff00000002000000020000;
		5'b00010:	xpb = 256'h000400000002000000020000000400000001fffffffe00000004000000040000;
		5'b00011:	xpb = 256'h000600000003000000030000000600000002fffffffd00000006000000060000;
		5'b00100:	xpb = 256'h000800000004000000040000000800000003fffffffc00000008000000080000;
		5'b00101:	xpb = 256'h000a00000005000000050000000a00000004fffffffb0000000a0000000a0000;
		5'b00110:	xpb = 256'h000c00000006000000060000000c00000005fffffffa0000000c0000000c0000;
		5'b00111:	xpb = 256'h000e00000007000000070000000e00000006fffffff90000000e0000000e0000;
		5'b01000:	xpb = 256'h001000000008000000080000001000000007fffffff800000010000000100000;
		5'b01001:	xpb = 256'h001200000009000000090000001200000008fffffff700000012000000120000;
		5'b01010:	xpb = 256'h00140000000a0000000a0000001400000009fffffff600000014000000140000;
		5'b01011:	xpb = 256'h00160000000b0000000b000000160000000afffffff500000016000000160000;
		5'b01100:	xpb = 256'h00180000000c0000000c000000180000000bfffffff400000018000000180000;
		5'b01101:	xpb = 256'h001a0000000d0000000d0000001a0000000cfffffff30000001a0000001a0000;
		5'b01110:	xpb = 256'h001c0000000e0000000e0000001c0000000dfffffff20000001c0000001c0000;
		5'b01111:	xpb = 256'h001e0000000f0000000f0000001e0000000efffffff10000001e0000001e0000;
		5'b10000:	xpb = 256'h00200000001000000010000000200000000ffffffff000000020000000200000;
		5'b10001:	xpb = 256'h002200000011000000110000002200000010ffffffef00000022000000220000;
		5'b10010:	xpb = 256'h002400000012000000120000002400000011ffffffee00000024000000240000;
		5'b10011:	xpb = 256'h002600000013000000130000002600000012ffffffed00000026000000260000;
		5'b10100:	xpb = 256'h002800000014000000140000002800000013ffffffec00000028000000280000;
		5'b10101:	xpb = 256'h002a00000015000000150000002a00000014ffffffeb0000002a0000002a0000;
		5'b10110:	xpb = 256'h002c00000016000000160000002c00000015ffffffea0000002c0000002c0000;
		5'b10111:	xpb = 256'h002e00000017000000170000002e00000016ffffffe90000002e0000002e0000;
		5'b11000:	xpb = 256'h003000000018000000180000003000000017ffffffe800000030000000300000;
		5'b11001:	xpb = 256'h003200000019000000190000003200000018ffffffe700000032000000320000;
		5'b11010:	xpb = 256'h00340000001a0000001a0000003400000019ffffffe600000034000000340000;
		5'b11011:	xpb = 256'h00360000001b0000001b000000360000001affffffe500000036000000360000;
		5'b11100:	xpb = 256'h00380000001c0000001c000000380000001bffffffe400000038000000380000;
		5'b11101:	xpb = 256'h003a0000001d0000001d0000003a0000001cffffffe30000003a0000003a0000;
		5'b11110:	xpb = 256'h003c0000001e0000001e0000003c0000001dffffffe20000003c0000003c0000;
		5'b11111:	xpb = 256'h003e0000001f0000001f0000003e0000001effffffe10000003e0000003e0000;
	endcase
end
endmodule

module xpb_29_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00400000002000000020000000400000001fffffffe000000040000000400000;
		6'b000010:	xpb = 256'h00800000004000000040000000800000003fffffffc000000080000000800000;
		6'b000011:	xpb = 256'h00c00000006000000060000000c00000005fffffffa0000000c0000000c00000;
		6'b000100:	xpb = 256'h01000000008000000080000001000000007fffffff8000000100000001000000;
		6'b000101:	xpb = 256'h0140000000a0000000a0000001400000009fffffff6000000140000001400000;
		6'b000110:	xpb = 256'h0180000000c0000000c000000180000000bfffffff4000000180000001800000;
		6'b000111:	xpb = 256'h01c0000000e0000000e0000001c0000000dfffffff20000001c0000001c00000;
		6'b001000:	xpb = 256'h0200000001000000010000000200000000ffffffff0000000200000002000000;
		6'b001001:	xpb = 256'h02400000012000000120000002400000011ffffffee000000240000002400000;
		6'b001010:	xpb = 256'h02800000014000000140000002800000013ffffffec000000280000002800000;
		6'b001011:	xpb = 256'h02c00000016000000160000002c00000015ffffffea0000002c0000002c00000;
		6'b001100:	xpb = 256'h03000000018000000180000003000000017ffffffe8000000300000003000000;
		6'b001101:	xpb = 256'h0340000001a0000001a0000003400000019ffffffe6000000340000003400000;
		6'b001110:	xpb = 256'h0380000001c0000001c000000380000001bffffffe4000000380000003800000;
		6'b001111:	xpb = 256'h03c0000001e0000001e0000003c0000001dffffffe20000003c0000003c00000;
		6'b010000:	xpb = 256'h0400000002000000020000000400000001fffffffe0000000400000004000000;
		6'b010001:	xpb = 256'h04400000022000000220000004400000021ffffffde000000440000004400000;
		6'b010010:	xpb = 256'h04800000024000000240000004800000023ffffffdc000000480000004800000;
		6'b010011:	xpb = 256'h04c00000026000000260000004c00000025ffffffda0000004c0000004c00000;
		6'b010100:	xpb = 256'h05000000028000000280000005000000027ffffffd8000000500000005000000;
		6'b010101:	xpb = 256'h0540000002a0000002a0000005400000029ffffffd6000000540000005400000;
		6'b010110:	xpb = 256'h0580000002c0000002c000000580000002bffffffd4000000580000005800000;
		6'b010111:	xpb = 256'h05c0000002e0000002e0000005c0000002dffffffd20000005c0000005c00000;
		6'b011000:	xpb = 256'h0600000003000000030000000600000002fffffffd0000000600000006000000;
		6'b011001:	xpb = 256'h06400000032000000320000006400000031ffffffce000000640000006400000;
		6'b011010:	xpb = 256'h06800000034000000340000006800000033ffffffcc000000680000006800000;
		6'b011011:	xpb = 256'h06c00000036000000360000006c00000035ffffffca0000006c0000006c00000;
		6'b011100:	xpb = 256'h07000000038000000380000007000000037ffffffc8000000700000007000000;
		6'b011101:	xpb = 256'h0740000003a0000003a0000007400000039ffffffc6000000740000007400000;
		6'b011110:	xpb = 256'h0780000003c0000003c000000780000003bffffffc4000000780000007800000;
		6'b011111:	xpb = 256'h07c0000003e0000003e0000007c0000003dffffffc20000007c0000007c00000;
		6'b100000:	xpb = 256'h0800000004000000040000000800000003fffffffc0000000800000008000000;
		6'b100001:	xpb = 256'h08400000042000000420000008400000041ffffffbe000000840000008400000;
		6'b100010:	xpb = 256'h08800000044000000440000008800000043ffffffbc000000880000008800000;
		6'b100011:	xpb = 256'h08c00000046000000460000008c00000045ffffffba0000008c0000008c00000;
		6'b100100:	xpb = 256'h09000000048000000480000009000000047ffffffb8000000900000009000000;
		6'b100101:	xpb = 256'h0940000004a0000004a0000009400000049ffffffb6000000940000009400000;
		6'b100110:	xpb = 256'h0980000004c0000004c000000980000004bffffffb4000000980000009800000;
		6'b100111:	xpb = 256'h09c0000004e0000004e0000009c0000004dffffffb20000009c0000009c00000;
		6'b101000:	xpb = 256'h0a00000005000000050000000a00000004fffffffb0000000a0000000a000000;
		6'b101001:	xpb = 256'h0a40000005200000052000000a400000051ffffffae000000a4000000a400000;
		6'b101010:	xpb = 256'h0a80000005400000054000000a800000053ffffffac000000a8000000a800000;
		6'b101011:	xpb = 256'h0ac0000005600000056000000ac00000055ffffffaa000000ac000000ac00000;
		6'b101100:	xpb = 256'h0b00000005800000058000000b000000057ffffffa8000000b0000000b000000;
		6'b101101:	xpb = 256'h0b40000005a0000005a000000b400000059ffffffa6000000b4000000b400000;
		6'b101110:	xpb = 256'h0b80000005c0000005c000000b80000005bffffffa4000000b8000000b800000;
		6'b101111:	xpb = 256'h0bc0000005e0000005e000000bc0000005dffffffa2000000bc000000bc00000;
		6'b110000:	xpb = 256'h0c00000006000000060000000c00000005fffffffa0000000c0000000c000000;
		6'b110001:	xpb = 256'h0c40000006200000062000000c400000061ffffff9e000000c4000000c400000;
		6'b110010:	xpb = 256'h0c80000006400000064000000c800000063ffffff9c000000c8000000c800000;
		6'b110011:	xpb = 256'h0cc0000006600000066000000cc00000065ffffff9a000000cc000000cc00000;
		6'b110100:	xpb = 256'h0d00000006800000068000000d000000067ffffff98000000d0000000d000000;
		6'b110101:	xpb = 256'h0d40000006a0000006a000000d400000069ffffff96000000d4000000d400000;
		6'b110110:	xpb = 256'h0d80000006c0000006c000000d80000006bffffff94000000d8000000d800000;
		6'b110111:	xpb = 256'h0dc0000006e0000006e000000dc0000006dffffff92000000dc000000dc00000;
		6'b111000:	xpb = 256'h0e00000007000000070000000e00000006fffffff90000000e0000000e000000;
		6'b111001:	xpb = 256'h0e40000007200000072000000e400000071ffffff8e000000e4000000e400000;
		6'b111010:	xpb = 256'h0e80000007400000074000000e800000073ffffff8c000000e8000000e800000;
		6'b111011:	xpb = 256'h0ec0000007600000076000000ec00000075ffffff8a000000ec000000ec00000;
		6'b111100:	xpb = 256'h0f00000007800000078000000f000000077ffffff88000000f0000000f000000;
		6'b111101:	xpb = 256'h0f40000007a0000007a000000f400000079ffffff86000000f4000000f400000;
		6'b111110:	xpb = 256'h0f80000007c0000007c000000f80000007bffffff84000000f8000000f800000;
		6'b111111:	xpb = 256'h0fc0000007e0000007e000000fc0000007dffffff82000000fc000000fc00000;
	endcase
end
endmodule

module xpb_29_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h1000000008000000080000001000000007fffffff80000001000000010000000;
		6'b000010:	xpb = 256'h200000001000000010000000200000000ffffffff00000002000000020000000;
		6'b000011:	xpb = 256'h3000000018000000180000003000000017ffffffe80000003000000030000000;
		6'b000100:	xpb = 256'h400000002000000020000000400000001fffffffe00000004000000040000000;
		6'b000101:	xpb = 256'h5000000028000000280000005000000027ffffffd80000005000000050000000;
		6'b000110:	xpb = 256'h600000003000000030000000600000002fffffffd00000006000000060000000;
		6'b000111:	xpb = 256'h7000000038000000380000007000000037ffffffc80000007000000070000000;
		6'b001000:	xpb = 256'h800000004000000040000000800000003fffffffc00000008000000080000000;
		6'b001001:	xpb = 256'h9000000048000000480000009000000047ffffffb80000009000000090000000;
		6'b001010:	xpb = 256'ha00000005000000050000000a00000004fffffffb0000000a0000000a0000000;
		6'b001011:	xpb = 256'hb00000005800000058000000b000000057ffffffa8000000b0000000b0000000;
		6'b001100:	xpb = 256'hc00000006000000060000000c00000005fffffffa0000000c0000000c0000000;
		6'b001101:	xpb = 256'hd00000006800000068000000d000000067ffffff98000000d0000000d0000000;
		6'b001110:	xpb = 256'he00000007000000070000000e00000006fffffff90000000e0000000e0000000;
		6'b001111:	xpb = 256'hf00000007800000078000000f000000077ffffff88000000f0000000f0000000;
		6'b010000:	xpb = 256'h0000000180000000800000010000000080000000800000000000000100000001;
		6'b010001:	xpb = 256'h1000000188000000880000011000000088000000780000001000000110000001;
		6'b010010:	xpb = 256'h2000000190000000900000012000000090000000700000002000000120000001;
		6'b010011:	xpb = 256'h3000000198000000980000013000000098000000680000003000000130000001;
		6'b010100:	xpb = 256'h40000001a0000000a000000140000000a0000000600000004000000140000001;
		6'b010101:	xpb = 256'h50000001a8000000a800000150000000a8000000580000005000000150000001;
		6'b010110:	xpb = 256'h60000001b0000000b000000160000000b0000000500000006000000160000001;
		6'b010111:	xpb = 256'h70000001b8000000b800000170000000b8000000480000007000000170000001;
		6'b011000:	xpb = 256'h80000001c0000000c000000180000000c0000000400000008000000180000001;
		6'b011001:	xpb = 256'h90000001c8000000c800000190000000c8000000380000009000000190000001;
		6'b011010:	xpb = 256'ha0000001d0000000d0000001a0000000d000000030000000a0000001a0000001;
		6'b011011:	xpb = 256'hb0000001d8000000d8000001b0000000d800000028000000b0000001b0000001;
		6'b011100:	xpb = 256'hc0000001e0000000e0000001c0000000e000000020000000c0000001c0000001;
		6'b011101:	xpb = 256'hd0000001e8000000e8000001d0000000e800000018000000d0000001d0000001;
		6'b011110:	xpb = 256'he0000001f0000000f0000001e0000000f000000010000000e0000001e0000001;
		6'b011111:	xpb = 256'hf0000001f8000000f8000001f0000000f800000008000000f0000001f0000001;
		6'b100000:	xpb = 256'h0000000300000001000000020000000100000001000000000000000200000002;
		6'b100001:	xpb = 256'h1000000308000001080000021000000108000000f80000001000000210000002;
		6'b100010:	xpb = 256'h2000000310000001100000022000000110000000f00000002000000220000002;
		6'b100011:	xpb = 256'h3000000318000001180000023000000118000000e80000003000000230000002;
		6'b100100:	xpb = 256'h4000000320000001200000024000000120000000e00000004000000240000002;
		6'b100101:	xpb = 256'h5000000328000001280000025000000128000000d80000005000000250000002;
		6'b100110:	xpb = 256'h6000000330000001300000026000000130000000d00000006000000260000002;
		6'b100111:	xpb = 256'h7000000338000001380000027000000138000000c80000007000000270000002;
		6'b101000:	xpb = 256'h8000000340000001400000028000000140000000c00000008000000280000002;
		6'b101001:	xpb = 256'h9000000348000001480000029000000148000000b80000009000000290000002;
		6'b101010:	xpb = 256'ha00000035000000150000002a000000150000000b0000000a0000002a0000002;
		6'b101011:	xpb = 256'hb00000035800000158000002b000000158000000a8000000b0000002b0000002;
		6'b101100:	xpb = 256'hc00000036000000160000002c000000160000000a0000000c0000002c0000002;
		6'b101101:	xpb = 256'hd00000036800000168000002d00000016800000098000000d0000002d0000002;
		6'b101110:	xpb = 256'he00000037000000170000002e00000017000000090000000e0000002e0000002;
		6'b101111:	xpb = 256'hf00000037800000178000002f00000017800000088000000f0000002f0000002;
		6'b110000:	xpb = 256'h0000000480000001800000030000000180000001800000000000000300000003;
		6'b110001:	xpb = 256'h1000000488000001880000031000000188000001780000001000000310000003;
		6'b110010:	xpb = 256'h2000000490000001900000032000000190000001700000002000000320000003;
		6'b110011:	xpb = 256'h3000000498000001980000033000000198000001680000003000000330000003;
		6'b110100:	xpb = 256'h40000004a0000001a000000340000001a0000001600000004000000340000003;
		6'b110101:	xpb = 256'h50000004a8000001a800000350000001a8000001580000005000000350000003;
		6'b110110:	xpb = 256'h60000004b0000001b000000360000001b0000001500000006000000360000003;
		6'b110111:	xpb = 256'h70000004b8000001b800000370000001b8000001480000007000000370000003;
		6'b111000:	xpb = 256'h80000004c0000001c000000380000001c0000001400000008000000380000003;
		6'b111001:	xpb = 256'h90000004c8000001c800000390000001c8000001380000009000000390000003;
		6'b111010:	xpb = 256'ha0000004d0000001d0000003a0000001d000000130000000a0000003a0000003;
		6'b111011:	xpb = 256'hb0000004d8000001d8000003b0000001d800000128000000b0000003b0000003;
		6'b111100:	xpb = 256'hc0000004e0000001e0000003c0000001e000000120000000c0000003c0000003;
		6'b111101:	xpb = 256'hd0000004e8000001e8000003d0000001e800000118000000d0000003d0000003;
		6'b111110:	xpb = 256'he0000004f0000001f0000003e0000001f000000110000000e0000003e0000003;
		6'b111111:	xpb = 256'hf0000004f8000001f8000003f0000001f800000108000000f0000003f0000003;
	endcase
end
endmodule

module xpb_30_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000300000001000000020000000100000001000000000000000200000002;
		5'b00010:	xpb = 256'h0000000600000002000000040000000200000002000000000000000400000004;
		5'b00011:	xpb = 256'h0000000900000003000000060000000300000003000000000000000600000006;
		5'b00100:	xpb = 256'h0000000c00000004000000080000000400000004000000000000000800000008;
		5'b00101:	xpb = 256'h0000000f000000050000000a0000000500000005000000000000000a0000000a;
		5'b00110:	xpb = 256'h00000012000000060000000c0000000600000006000000000000000c0000000c;
		5'b00111:	xpb = 256'h00000015000000070000000e0000000700000007000000000000000e0000000e;
		5'b01000:	xpb = 256'h0000001800000008000000100000000800000008000000000000001000000010;
		5'b01001:	xpb = 256'h0000001b00000009000000120000000900000009000000000000001200000012;
		5'b01010:	xpb = 256'h0000001e0000000a000000140000000a0000000a000000000000001400000014;
		5'b01011:	xpb = 256'h000000210000000b000000160000000b0000000b000000000000001600000016;
		5'b01100:	xpb = 256'h000000240000000c000000180000000c0000000c000000000000001800000018;
		5'b01101:	xpb = 256'h000000270000000d0000001a0000000d0000000d000000000000001a0000001a;
		5'b01110:	xpb = 256'h0000002a0000000e0000001c0000000e0000000e000000000000001c0000001c;
		5'b01111:	xpb = 256'h0000002d0000000f0000001e0000000f0000000f000000000000001e0000001e;
		5'b10000:	xpb = 256'h0000003000000010000000200000001000000010000000000000002000000020;
		5'b10001:	xpb = 256'h0000003300000011000000220000001100000011000000000000002200000022;
		5'b10010:	xpb = 256'h0000003600000012000000240000001200000012000000000000002400000024;
		5'b10011:	xpb = 256'h0000003900000013000000260000001300000013000000000000002600000026;
		5'b10100:	xpb = 256'h0000003c00000014000000280000001400000014000000000000002800000028;
		5'b10101:	xpb = 256'h0000003f000000150000002a0000001500000015000000000000002a0000002a;
		5'b10110:	xpb = 256'h00000042000000160000002c0000001600000016000000000000002c0000002c;
		5'b10111:	xpb = 256'h00000045000000170000002e0000001700000017000000000000002e0000002e;
		5'b11000:	xpb = 256'h0000004800000018000000300000001800000018000000000000003000000030;
		5'b11001:	xpb = 256'h0000004b00000019000000320000001900000019000000000000003200000032;
		5'b11010:	xpb = 256'h0000004e0000001a000000340000001a0000001a000000000000003400000034;
		5'b11011:	xpb = 256'h000000510000001b000000360000001b0000001b000000000000003600000036;
		5'b11100:	xpb = 256'h000000540000001c000000380000001c0000001c000000000000003800000038;
		5'b11101:	xpb = 256'h000000570000001d0000003a0000001d0000001d000000000000003a0000003a;
		5'b11110:	xpb = 256'h0000005a0000001e0000003c0000001e0000001e000000000000003c0000003c;
		5'b11111:	xpb = 256'h0000005d0000001f0000003e0000001f0000001f000000000000003e0000003e;
	endcase
end
endmodule

module xpb_30_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000006000000020000000400000002000000020000000000000004000000040;
		6'b000010:	xpb = 256'h000000c000000040000000800000004000000040000000000000008000000080;
		6'b000011:	xpb = 256'h0000012000000060000000c0000000600000006000000000000000c0000000c0;
		6'b000100:	xpb = 256'h0000018000000080000001000000008000000080000000000000010000000100;
		6'b000101:	xpb = 256'h000001e0000000a000000140000000a0000000a0000000000000014000000140;
		6'b000110:	xpb = 256'h00000240000000c000000180000000c0000000c0000000000000018000000180;
		6'b000111:	xpb = 256'h000002a0000000e0000001c0000000e0000000e000000000000001c0000001c0;
		6'b001000:	xpb = 256'h0000030000000100000002000000010000000100000000000000020000000200;
		6'b001001:	xpb = 256'h0000036000000120000002400000012000000120000000000000024000000240;
		6'b001010:	xpb = 256'h000003c000000140000002800000014000000140000000000000028000000280;
		6'b001011:	xpb = 256'h0000042000000160000002c0000001600000016000000000000002c0000002c0;
		6'b001100:	xpb = 256'h0000048000000180000003000000018000000180000000000000030000000300;
		6'b001101:	xpb = 256'h000004e0000001a000000340000001a0000001a0000000000000034000000340;
		6'b001110:	xpb = 256'h00000540000001c000000380000001c0000001c0000000000000038000000380;
		6'b001111:	xpb = 256'h000005a0000001e0000003c0000001e0000001e000000000000003c0000003c0;
		6'b010000:	xpb = 256'h0000060000000200000004000000020000000200000000000000040000000400;
		6'b010001:	xpb = 256'h0000066000000220000004400000022000000220000000000000044000000440;
		6'b010010:	xpb = 256'h000006c000000240000004800000024000000240000000000000048000000480;
		6'b010011:	xpb = 256'h0000072000000260000004c0000002600000026000000000000004c0000004c0;
		6'b010100:	xpb = 256'h0000078000000280000005000000028000000280000000000000050000000500;
		6'b010101:	xpb = 256'h000007e0000002a000000540000002a0000002a0000000000000054000000540;
		6'b010110:	xpb = 256'h00000840000002c000000580000002c0000002c0000000000000058000000580;
		6'b010111:	xpb = 256'h000008a0000002e0000005c0000002e0000002e000000000000005c0000005c0;
		6'b011000:	xpb = 256'h0000090000000300000006000000030000000300000000000000060000000600;
		6'b011001:	xpb = 256'h0000096000000320000006400000032000000320000000000000064000000640;
		6'b011010:	xpb = 256'h000009c000000340000006800000034000000340000000000000068000000680;
		6'b011011:	xpb = 256'h00000a2000000360000006c0000003600000036000000000000006c0000006c0;
		6'b011100:	xpb = 256'h00000a8000000380000007000000038000000380000000000000070000000700;
		6'b011101:	xpb = 256'h00000ae0000003a000000740000003a0000003a0000000000000074000000740;
		6'b011110:	xpb = 256'h00000b40000003c000000780000003c0000003c0000000000000078000000780;
		6'b011111:	xpb = 256'h00000ba0000003e0000007c0000003e0000003e000000000000007c0000007c0;
		6'b100000:	xpb = 256'h00000c0000000400000008000000040000000400000000000000080000000800;
		6'b100001:	xpb = 256'h00000c6000000420000008400000042000000420000000000000084000000840;
		6'b100010:	xpb = 256'h00000cc000000440000008800000044000000440000000000000088000000880;
		6'b100011:	xpb = 256'h00000d2000000460000008c0000004600000046000000000000008c0000008c0;
		6'b100100:	xpb = 256'h00000d8000000480000009000000048000000480000000000000090000000900;
		6'b100101:	xpb = 256'h00000de0000004a000000940000004a0000004a0000000000000094000000940;
		6'b100110:	xpb = 256'h00000e40000004c000000980000004c0000004c0000000000000098000000980;
		6'b100111:	xpb = 256'h00000ea0000004e0000009c0000004e0000004e000000000000009c0000009c0;
		6'b101000:	xpb = 256'h00000f000000050000000a0000000500000005000000000000000a0000000a00;
		6'b101001:	xpb = 256'h00000f600000052000000a4000000520000005200000000000000a4000000a40;
		6'b101010:	xpb = 256'h00000fc00000054000000a8000000540000005400000000000000a8000000a80;
		6'b101011:	xpb = 256'h000010200000056000000ac000000560000005600000000000000ac000000ac0;
		6'b101100:	xpb = 256'h000010800000058000000b0000000580000005800000000000000b0000000b00;
		6'b101101:	xpb = 256'h000010e0000005a000000b40000005a0000005a00000000000000b4000000b40;
		6'b101110:	xpb = 256'h00001140000005c000000b80000005c0000005c00000000000000b8000000b80;
		6'b101111:	xpb = 256'h000011a0000005e000000bc0000005e0000005e00000000000000bc000000bc0;
		6'b110000:	xpb = 256'h000012000000060000000c0000000600000006000000000000000c0000000c00;
		6'b110001:	xpb = 256'h000012600000062000000c4000000620000006200000000000000c4000000c40;
		6'b110010:	xpb = 256'h000012c00000064000000c8000000640000006400000000000000c8000000c80;
		6'b110011:	xpb = 256'h000013200000066000000cc000000660000006600000000000000cc000000cc0;
		6'b110100:	xpb = 256'h000013800000068000000d0000000680000006800000000000000d0000000d00;
		6'b110101:	xpb = 256'h000013e0000006a000000d40000006a0000006a00000000000000d4000000d40;
		6'b110110:	xpb = 256'h00001440000006c000000d80000006c0000006c00000000000000d8000000d80;
		6'b110111:	xpb = 256'h000014a0000006e000000dc0000006e0000006e00000000000000dc000000dc0;
		6'b111000:	xpb = 256'h000015000000070000000e0000000700000007000000000000000e0000000e00;
		6'b111001:	xpb = 256'h000015600000072000000e4000000720000007200000000000000e4000000e40;
		6'b111010:	xpb = 256'h000015c00000074000000e8000000740000007400000000000000e8000000e80;
		6'b111011:	xpb = 256'h000016200000076000000ec000000760000007600000000000000ec000000ec0;
		6'b111100:	xpb = 256'h000016800000078000000f0000000780000007800000000000000f0000000f00;
		6'b111101:	xpb = 256'h000016e0000007a000000f40000007a0000007a00000000000000f4000000f40;
		6'b111110:	xpb = 256'h00001740000007c000000f80000007c0000007c00000000000000f8000000f80;
		6'b111111:	xpb = 256'h000017a0000007e000000fc0000007e0000007e00000000000000fc000000fc0;
	endcase
end
endmodule

module xpb_30_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000180000000800000010000000080000000800000000000000100000001000;
		6'b000010:	xpb = 256'h0000300000001000000020000000100000001000000000000000200000002000;
		6'b000011:	xpb = 256'h0000480000001800000030000000180000001800000000000000300000003000;
		6'b000100:	xpb = 256'h0000600000002000000040000000200000002000000000000000400000004000;
		6'b000101:	xpb = 256'h0000780000002800000050000000280000002800000000000000500000005000;
		6'b000110:	xpb = 256'h0000900000003000000060000000300000003000000000000000600000006000;
		6'b000111:	xpb = 256'h0000a80000003800000070000000380000003800000000000000700000007000;
		6'b001000:	xpb = 256'h0000c00000004000000080000000400000004000000000000000800000008000;
		6'b001001:	xpb = 256'h0000d80000004800000090000000480000004800000000000000900000009000;
		6'b001010:	xpb = 256'h0000f000000050000000a0000000500000005000000000000000a0000000a000;
		6'b001011:	xpb = 256'h00010800000058000000b0000000580000005800000000000000b0000000b000;
		6'b001100:	xpb = 256'h00012000000060000000c0000000600000006000000000000000c0000000c000;
		6'b001101:	xpb = 256'h00013800000068000000d0000000680000006800000000000000d0000000d000;
		6'b001110:	xpb = 256'h00015000000070000000e0000000700000007000000000000000e0000000e000;
		6'b001111:	xpb = 256'h00016800000078000000f0000000780000007800000000000000f0000000f000;
		6'b010000:	xpb = 256'h0001800000008000000100000000800000008000000000000001000000010000;
		6'b010001:	xpb = 256'h0001980000008800000110000000880000008800000000000001100000011000;
		6'b010010:	xpb = 256'h0001b00000009000000120000000900000009000000000000001200000012000;
		6'b010011:	xpb = 256'h0001c80000009800000130000000980000009800000000000001300000013000;
		6'b010100:	xpb = 256'h0001e0000000a000000140000000a0000000a000000000000001400000014000;
		6'b010101:	xpb = 256'h0001f8000000a800000150000000a8000000a800000000000001500000015000;
		6'b010110:	xpb = 256'h000210000000b000000160000000b0000000b000000000000001600000016000;
		6'b010111:	xpb = 256'h000228000000b800000170000000b8000000b800000000000001700000017000;
		6'b011000:	xpb = 256'h000240000000c000000180000000c0000000c000000000000001800000018000;
		6'b011001:	xpb = 256'h000258000000c800000190000000c8000000c800000000000001900000019000;
		6'b011010:	xpb = 256'h000270000000d0000001a0000000d0000000d000000000000001a0000001a000;
		6'b011011:	xpb = 256'h000288000000d8000001b0000000d8000000d800000000000001b0000001b000;
		6'b011100:	xpb = 256'h0002a0000000e0000001c0000000e0000000e000000000000001c0000001c000;
		6'b011101:	xpb = 256'h0002b8000000e8000001d0000000e8000000e800000000000001d0000001d000;
		6'b011110:	xpb = 256'h0002d0000000f0000001e0000000f0000000f000000000000001e0000001e000;
		6'b011111:	xpb = 256'h0002e8000000f8000001f0000000f8000000f800000000000001f0000001f000;
		6'b100000:	xpb = 256'h0003000000010000000200000001000000010000000000000002000000020000;
		6'b100001:	xpb = 256'h0003180000010800000210000001080000010800000000000002100000021000;
		6'b100010:	xpb = 256'h0003300000011000000220000001100000011000000000000002200000022000;
		6'b100011:	xpb = 256'h0003480000011800000230000001180000011800000000000002300000023000;
		6'b100100:	xpb = 256'h0003600000012000000240000001200000012000000000000002400000024000;
		6'b100101:	xpb = 256'h0003780000012800000250000001280000012800000000000002500000025000;
		6'b100110:	xpb = 256'h0003900000013000000260000001300000013000000000000002600000026000;
		6'b100111:	xpb = 256'h0003a80000013800000270000001380000013800000000000002700000027000;
		6'b101000:	xpb = 256'h0003c00000014000000280000001400000014000000000000002800000028000;
		6'b101001:	xpb = 256'h0003d80000014800000290000001480000014800000000000002900000029000;
		6'b101010:	xpb = 256'h0003f000000150000002a0000001500000015000000000000002a0000002a000;
		6'b101011:	xpb = 256'h00040800000158000002b0000001580000015800000000000002b0000002b000;
		6'b101100:	xpb = 256'h00042000000160000002c0000001600000016000000000000002c0000002c000;
		6'b101101:	xpb = 256'h00043800000168000002d0000001680000016800000000000002d0000002d000;
		6'b101110:	xpb = 256'h00045000000170000002e0000001700000017000000000000002e0000002e000;
		6'b101111:	xpb = 256'h00046800000178000002f0000001780000017800000000000002f0000002f000;
		6'b110000:	xpb = 256'h0004800000018000000300000001800000018000000000000003000000030000;
		6'b110001:	xpb = 256'h0004980000018800000310000001880000018800000000000003100000031000;
		6'b110010:	xpb = 256'h0004b00000019000000320000001900000019000000000000003200000032000;
		6'b110011:	xpb = 256'h0004c80000019800000330000001980000019800000000000003300000033000;
		6'b110100:	xpb = 256'h0004e0000001a000000340000001a0000001a000000000000003400000034000;
		6'b110101:	xpb = 256'h0004f8000001a800000350000001a8000001a800000000000003500000035000;
		6'b110110:	xpb = 256'h000510000001b000000360000001b0000001b000000000000003600000036000;
		6'b110111:	xpb = 256'h000528000001b800000370000001b8000001b800000000000003700000037000;
		6'b111000:	xpb = 256'h000540000001c000000380000001c0000001c000000000000003800000038000;
		6'b111001:	xpb = 256'h000558000001c800000390000001c8000001c800000000000003900000039000;
		6'b111010:	xpb = 256'h000570000001d0000003a0000001d0000001d000000000000003a0000003a000;
		6'b111011:	xpb = 256'h000588000001d8000003b0000001d8000001d800000000000003b0000003b000;
		6'b111100:	xpb = 256'h0005a0000001e0000003c0000001e0000001e000000000000003c0000003c000;
		6'b111101:	xpb = 256'h0005b8000001e8000003d0000001e8000001e800000000000003d0000003d000;
		6'b111110:	xpb = 256'h0005d0000001f0000003e0000001f0000001f000000000000003e0000003e000;
		6'b111111:	xpb = 256'h0005e8000001f8000003f0000001f8000001f800000000000003f0000003f000;
	endcase
end
endmodule

module xpb_31_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0003000000010000000200000001000000010000000000000002000000020000;
		5'b00010:	xpb = 256'h0006000000020000000400000002000000020000000000000004000000040000;
		5'b00011:	xpb = 256'h0009000000030000000600000003000000030000000000000006000000060000;
		5'b00100:	xpb = 256'h000c000000040000000800000004000000040000000000000008000000080000;
		5'b00101:	xpb = 256'h000f000000050000000a0000000500000005000000000000000a0000000a0000;
		5'b00110:	xpb = 256'h0012000000060000000c0000000600000006000000000000000c0000000c0000;
		5'b00111:	xpb = 256'h0015000000070000000e0000000700000007000000000000000e0000000e0000;
		5'b01000:	xpb = 256'h0018000000080000001000000008000000080000000000000010000000100000;
		5'b01001:	xpb = 256'h001b000000090000001200000009000000090000000000000012000000120000;
		5'b01010:	xpb = 256'h001e0000000a000000140000000a0000000a0000000000000014000000140000;
		5'b01011:	xpb = 256'h00210000000b000000160000000b0000000b0000000000000016000000160000;
		5'b01100:	xpb = 256'h00240000000c000000180000000c0000000c0000000000000018000000180000;
		5'b01101:	xpb = 256'h00270000000d0000001a0000000d0000000d000000000000001a0000001a0000;
		5'b01110:	xpb = 256'h002a0000000e0000001c0000000e0000000e000000000000001c0000001c0000;
		5'b01111:	xpb = 256'h002d0000000f0000001e0000000f0000000f000000000000001e0000001e0000;
		5'b10000:	xpb = 256'h0030000000100000002000000010000000100000000000000020000000200000;
		5'b10001:	xpb = 256'h0033000000110000002200000011000000110000000000000022000000220000;
		5'b10010:	xpb = 256'h0036000000120000002400000012000000120000000000000024000000240000;
		5'b10011:	xpb = 256'h0039000000130000002600000013000000130000000000000026000000260000;
		5'b10100:	xpb = 256'h003c000000140000002800000014000000140000000000000028000000280000;
		5'b10101:	xpb = 256'h003f000000150000002a0000001500000015000000000000002a0000002a0000;
		5'b10110:	xpb = 256'h0042000000160000002c0000001600000016000000000000002c0000002c0000;
		5'b10111:	xpb = 256'h0045000000170000002e0000001700000017000000000000002e0000002e0000;
		5'b11000:	xpb = 256'h0048000000180000003000000018000000180000000000000030000000300000;
		5'b11001:	xpb = 256'h004b000000190000003200000019000000190000000000000032000000320000;
		5'b11010:	xpb = 256'h004e0000001a000000340000001a0000001a0000000000000034000000340000;
		5'b11011:	xpb = 256'h00510000001b000000360000001b0000001b0000000000000036000000360000;
		5'b11100:	xpb = 256'h00540000001c000000380000001c0000001c0000000000000038000000380000;
		5'b11101:	xpb = 256'h00570000001d0000003a0000001d0000001d000000000000003a0000003a0000;
		5'b11110:	xpb = 256'h005a0000001e0000003c0000001e0000001e000000000000003c0000003c0000;
		5'b11111:	xpb = 256'h005d0000001f0000003e0000001f0000001f000000000000003e0000003e0000;
	endcase
end
endmodule

module xpb_31_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0060000000200000004000000020000000200000000000000040000000400000;
		6'b000010:	xpb = 256'h00c0000000400000008000000040000000400000000000000080000000800000;
		6'b000011:	xpb = 256'h012000000060000000c0000000600000006000000000000000c0000000c00000;
		6'b000100:	xpb = 256'h0180000000800000010000000080000000800000000000000100000001000000;
		6'b000101:	xpb = 256'h01e0000000a000000140000000a0000000a00000000000000140000001400000;
		6'b000110:	xpb = 256'h0240000000c000000180000000c0000000c00000000000000180000001800000;
		6'b000111:	xpb = 256'h02a0000000e0000001c0000000e0000000e000000000000001c0000001c00000;
		6'b001000:	xpb = 256'h0300000001000000020000000100000001000000000000000200000002000000;
		6'b001001:	xpb = 256'h0360000001200000024000000120000001200000000000000240000002400000;
		6'b001010:	xpb = 256'h03c0000001400000028000000140000001400000000000000280000002800000;
		6'b001011:	xpb = 256'h042000000160000002c0000001600000016000000000000002c0000002c00000;
		6'b001100:	xpb = 256'h0480000001800000030000000180000001800000000000000300000003000000;
		6'b001101:	xpb = 256'h04e0000001a000000340000001a0000001a00000000000000340000003400000;
		6'b001110:	xpb = 256'h0540000001c000000380000001c0000001c00000000000000380000003800000;
		6'b001111:	xpb = 256'h05a0000001e0000003c0000001e0000001e000000000000003c0000003c00000;
		6'b010000:	xpb = 256'h0600000002000000040000000200000002000000000000000400000004000000;
		6'b010001:	xpb = 256'h0660000002200000044000000220000002200000000000000440000004400000;
		6'b010010:	xpb = 256'h06c0000002400000048000000240000002400000000000000480000004800000;
		6'b010011:	xpb = 256'h072000000260000004c0000002600000026000000000000004c0000004c00000;
		6'b010100:	xpb = 256'h0780000002800000050000000280000002800000000000000500000005000000;
		6'b010101:	xpb = 256'h07e0000002a000000540000002a0000002a00000000000000540000005400000;
		6'b010110:	xpb = 256'h0840000002c000000580000002c0000002c00000000000000580000005800000;
		6'b010111:	xpb = 256'h08a0000002e0000005c0000002e0000002e000000000000005c0000005c00000;
		6'b011000:	xpb = 256'h0900000003000000060000000300000003000000000000000600000006000000;
		6'b011001:	xpb = 256'h0960000003200000064000000320000003200000000000000640000006400000;
		6'b011010:	xpb = 256'h09c0000003400000068000000340000003400000000000000680000006800000;
		6'b011011:	xpb = 256'h0a2000000360000006c0000003600000036000000000000006c0000006c00000;
		6'b011100:	xpb = 256'h0a80000003800000070000000380000003800000000000000700000007000000;
		6'b011101:	xpb = 256'h0ae0000003a000000740000003a0000003a00000000000000740000007400000;
		6'b011110:	xpb = 256'h0b40000003c000000780000003c0000003c00000000000000780000007800000;
		6'b011111:	xpb = 256'h0ba0000003e0000007c0000003e0000003e000000000000007c0000007c00000;
		6'b100000:	xpb = 256'h0c00000004000000080000000400000004000000000000000800000008000000;
		6'b100001:	xpb = 256'h0c60000004200000084000000420000004200000000000000840000008400000;
		6'b100010:	xpb = 256'h0cc0000004400000088000000440000004400000000000000880000008800000;
		6'b100011:	xpb = 256'h0d2000000460000008c0000004600000046000000000000008c0000008c00000;
		6'b100100:	xpb = 256'h0d80000004800000090000000480000004800000000000000900000009000000;
		6'b100101:	xpb = 256'h0de0000004a000000940000004a0000004a00000000000000940000009400000;
		6'b100110:	xpb = 256'h0e40000004c000000980000004c0000004c00000000000000980000009800000;
		6'b100111:	xpb = 256'h0ea0000004e0000009c0000004e0000004e000000000000009c0000009c00000;
		6'b101000:	xpb = 256'h0f000000050000000a0000000500000005000000000000000a0000000a000000;
		6'b101001:	xpb = 256'h0f600000052000000a4000000520000005200000000000000a4000000a400000;
		6'b101010:	xpb = 256'h0fc00000054000000a8000000540000005400000000000000a8000000a800000;
		6'b101011:	xpb = 256'h10200000056000000ac000000560000005600000000000000ac000000ac00000;
		6'b101100:	xpb = 256'h10800000058000000b0000000580000005800000000000000b0000000b000000;
		6'b101101:	xpb = 256'h10e0000005a000000b40000005a0000005a00000000000000b4000000b400000;
		6'b101110:	xpb = 256'h1140000005c000000b80000005c0000005c00000000000000b8000000b800000;
		6'b101111:	xpb = 256'h11a0000005e000000bc0000005e0000005e00000000000000bc000000bc00000;
		6'b110000:	xpb = 256'h12000000060000000c0000000600000006000000000000000c0000000c000000;
		6'b110001:	xpb = 256'h12600000062000000c4000000620000006200000000000000c4000000c400000;
		6'b110010:	xpb = 256'h12c00000064000000c8000000640000006400000000000000c8000000c800000;
		6'b110011:	xpb = 256'h13200000066000000cc000000660000006600000000000000cc000000cc00000;
		6'b110100:	xpb = 256'h13800000068000000d0000000680000006800000000000000d0000000d000000;
		6'b110101:	xpb = 256'h13e0000006a000000d40000006a0000006a00000000000000d4000000d400000;
		6'b110110:	xpb = 256'h1440000006c000000d80000006c0000006c00000000000000d8000000d800000;
		6'b110111:	xpb = 256'h14a0000006e000000dc0000006e0000006e00000000000000dc000000dc00000;
		6'b111000:	xpb = 256'h15000000070000000e0000000700000007000000000000000e0000000e000000;
		6'b111001:	xpb = 256'h15600000072000000e4000000720000007200000000000000e4000000e400000;
		6'b111010:	xpb = 256'h15c00000074000000e8000000740000007400000000000000e8000000e800000;
		6'b111011:	xpb = 256'h16200000076000000ec000000760000007600000000000000ec000000ec00000;
		6'b111100:	xpb = 256'h16800000078000000f0000000780000007800000000000000f0000000f000000;
		6'b111101:	xpb = 256'h16e0000007a000000f40000007a0000007a00000000000000f4000000f400000;
		6'b111110:	xpb = 256'h1740000007c000000f80000007c0000007c00000000000000f8000000f800000;
		6'b111111:	xpb = 256'h17a0000007e000000fc0000007e0000007e00000000000000fc000000fc00000;
	endcase
end
endmodule

module xpb_31_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h1800000008000000100000000800000008000000000000001000000010000000;
		6'b000010:	xpb = 256'h3000000010000000200000001000000010000000000000002000000020000000;
		6'b000011:	xpb = 256'h4800000018000000300000001800000018000000000000003000000030000000;
		6'b000100:	xpb = 256'h6000000020000000400000002000000020000000000000004000000040000000;
		6'b000101:	xpb = 256'h7800000028000000500000002800000028000000000000005000000050000000;
		6'b000110:	xpb = 256'h9000000030000000600000003000000030000000000000006000000060000000;
		6'b000111:	xpb = 256'ha800000038000000700000003800000038000000000000007000000070000000;
		6'b001000:	xpb = 256'hc000000040000000800000004000000040000000000000008000000080000000;
		6'b001001:	xpb = 256'hd800000048000000900000004800000048000000000000009000000090000000;
		6'b001010:	xpb = 256'hf000000050000000a0000000500000005000000000000000a0000000a0000000;
		6'b001011:	xpb = 256'h0800000158000000b00000005800000058000000ffffffffb0000000b0000001;
		6'b001100:	xpb = 256'h2000000160000000c00000006000000060000000ffffffffc0000000c0000001;
		6'b001101:	xpb = 256'h3800000168000000d00000006800000068000000ffffffffd0000000d0000001;
		6'b001110:	xpb = 256'h5000000170000000e00000007000000070000000ffffffffe0000000e0000001;
		6'b001111:	xpb = 256'h6800000178000000f00000007800000078000000fffffffff0000000f0000001;
		6'b010000:	xpb = 256'h8000000180000001000000008000000080000001000000000000000100000001;
		6'b010001:	xpb = 256'h9800000188000001100000008800000088000001000000001000000110000001;
		6'b010010:	xpb = 256'hb000000190000001200000009000000090000001000000002000000120000001;
		6'b010011:	xpb = 256'hc800000198000001300000009800000098000001000000003000000130000001;
		6'b010100:	xpb = 256'he0000001a000000140000000a0000000a0000001000000004000000140000001;
		6'b010101:	xpb = 256'hf8000001a800000150000000a8000000a8000001000000005000000150000001;
		6'b010110:	xpb = 256'h10000002b000000160000000b0000000b0000001ffffffff6000000160000002;
		6'b010111:	xpb = 256'h28000002b800000170000000b8000000b8000001ffffffff7000000170000002;
		6'b011000:	xpb = 256'h40000002c000000180000000c0000000c0000001ffffffff8000000180000002;
		6'b011001:	xpb = 256'h58000002c800000190000000c8000000c8000001ffffffff9000000190000002;
		6'b011010:	xpb = 256'h70000002d0000001a0000000d0000000d0000001ffffffffa0000001a0000002;
		6'b011011:	xpb = 256'h88000002d8000001b0000000d8000000d8000001ffffffffb0000001b0000002;
		6'b011100:	xpb = 256'ha0000002e0000001c0000000e0000000e0000001ffffffffc0000001c0000002;
		6'b011101:	xpb = 256'hb8000002e8000001d0000000e8000000e8000001ffffffffd0000001d0000002;
		6'b011110:	xpb = 256'hd0000002f0000001e0000000f0000000f0000001ffffffffe0000001e0000002;
		6'b011111:	xpb = 256'he8000002f8000001f0000000f8000000f8000001fffffffff0000001f0000002;
		6'b100000:	xpb = 256'h0000000400000002000000010000000100000002ffffffff0000000200000003;
		6'b100001:	xpb = 256'h1800000408000002100000010800000108000002ffffffff1000000210000003;
		6'b100010:	xpb = 256'h3000000410000002200000011000000110000002ffffffff2000000220000003;
		6'b100011:	xpb = 256'h4800000418000002300000011800000118000002ffffffff3000000230000003;
		6'b100100:	xpb = 256'h6000000420000002400000012000000120000002ffffffff4000000240000003;
		6'b100101:	xpb = 256'h7800000428000002500000012800000128000002ffffffff5000000250000003;
		6'b100110:	xpb = 256'h9000000430000002600000013000000130000002ffffffff6000000260000003;
		6'b100111:	xpb = 256'ha800000438000002700000013800000138000002ffffffff7000000270000003;
		6'b101000:	xpb = 256'hc000000440000002800000014000000140000002ffffffff8000000280000003;
		6'b101001:	xpb = 256'hd800000448000002900000014800000148000002ffffffff9000000290000003;
		6'b101010:	xpb = 256'hf000000450000002a00000015000000150000002ffffffffa0000002a0000003;
		6'b101011:	xpb = 256'h0800000558000002b00000015800000158000003fffffffeb0000002b0000004;
		6'b101100:	xpb = 256'h2000000560000002c00000016000000160000003fffffffec0000002c0000004;
		6'b101101:	xpb = 256'h3800000568000002d00000016800000168000003fffffffed0000002d0000004;
		6'b101110:	xpb = 256'h5000000570000002e00000017000000170000003fffffffee0000002e0000004;
		6'b101111:	xpb = 256'h6800000578000002f00000017800000178000003fffffffef0000002f0000004;
		6'b110000:	xpb = 256'h8000000580000003000000018000000180000003ffffffff0000000300000004;
		6'b110001:	xpb = 256'h9800000588000003100000018800000188000003ffffffff1000000310000004;
		6'b110010:	xpb = 256'hb000000590000003200000019000000190000003ffffffff2000000320000004;
		6'b110011:	xpb = 256'hc800000598000003300000019800000198000003ffffffff3000000330000004;
		6'b110100:	xpb = 256'he0000005a000000340000001a0000001a0000003ffffffff4000000340000004;
		6'b110101:	xpb = 256'hf8000005a800000350000001a8000001a8000003ffffffff5000000350000004;
		6'b110110:	xpb = 256'h10000006b000000360000001b0000001b0000004fffffffe6000000360000005;
		6'b110111:	xpb = 256'h28000006b800000370000001b8000001b8000004fffffffe7000000370000005;
		6'b111000:	xpb = 256'h40000006c000000380000001c0000001c0000004fffffffe8000000380000005;
		6'b111001:	xpb = 256'h58000006c800000390000001c8000001c8000004fffffffe9000000390000005;
		6'b111010:	xpb = 256'h70000006d0000003a0000001d0000001d0000004fffffffea0000003a0000005;
		6'b111011:	xpb = 256'h88000006d8000003b0000001d8000001d8000004fffffffeb0000003b0000005;
		6'b111100:	xpb = 256'ha0000006e0000003c0000001e0000001e0000004fffffffec0000003c0000005;
		6'b111101:	xpb = 256'hb8000006e8000003d0000001e8000001e8000004fffffffed0000003d0000005;
		6'b111110:	xpb = 256'hd0000006f0000003e0000001f0000001f0000004fffffffee0000003e0000005;
		6'b111111:	xpb = 256'he8000006f8000003f0000001f8000001f8000004fffffffef0000003f0000005;
	endcase
end
endmodule

module xpb_32_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000400000002000000010000000100000002ffffffff0000000200000003;
		5'b00010:	xpb = 256'h0000000800000004000000020000000200000005fffffffe0000000400000006;
		5'b00011:	xpb = 256'h0000000c00000006000000030000000300000008fffffffd0000000600000009;
		5'b00100:	xpb = 256'h000000100000000800000004000000040000000bfffffffc000000080000000c;
		5'b00101:	xpb = 256'h000000140000000a00000005000000050000000efffffffb0000000a0000000f;
		5'b00110:	xpb = 256'h000000180000000c000000060000000600000011fffffffa0000000c00000012;
		5'b00111:	xpb = 256'h0000001c0000000e000000070000000700000014fffffff90000000e00000015;
		5'b01000:	xpb = 256'h0000002000000010000000080000000800000017fffffff80000001000000018;
		5'b01001:	xpb = 256'h000000240000001200000009000000090000001afffffff7000000120000001b;
		5'b01010:	xpb = 256'h00000028000000140000000a0000000a0000001dfffffff6000000140000001e;
		5'b01011:	xpb = 256'h0000002c000000160000000b0000000b00000020fffffff50000001600000021;
		5'b01100:	xpb = 256'h00000030000000180000000c0000000c00000023fffffff40000001800000024;
		5'b01101:	xpb = 256'h000000340000001a0000000d0000000d00000026fffffff30000001a00000027;
		5'b01110:	xpb = 256'h000000380000001c0000000e0000000e00000029fffffff20000001c0000002a;
		5'b01111:	xpb = 256'h0000003c0000001e0000000f0000000f0000002cfffffff10000001e0000002d;
		5'b10000:	xpb = 256'h000000400000002000000010000000100000002ffffffff00000002000000030;
		5'b10001:	xpb = 256'h0000004400000022000000110000001100000032ffffffef0000002200000033;
		5'b10010:	xpb = 256'h0000004800000024000000120000001200000035ffffffee0000002400000036;
		5'b10011:	xpb = 256'h0000004c00000026000000130000001300000038ffffffed0000002600000039;
		5'b10100:	xpb = 256'h000000500000002800000014000000140000003bffffffec000000280000003c;
		5'b10101:	xpb = 256'h000000540000002a00000015000000150000003effffffeb0000002a0000003f;
		5'b10110:	xpb = 256'h000000580000002c000000160000001600000041ffffffea0000002c00000042;
		5'b10111:	xpb = 256'h0000005c0000002e000000170000001700000044ffffffe90000002e00000045;
		5'b11000:	xpb = 256'h0000006000000030000000180000001800000047ffffffe80000003000000048;
		5'b11001:	xpb = 256'h000000640000003200000019000000190000004affffffe7000000320000004b;
		5'b11010:	xpb = 256'h00000068000000340000001a0000001a0000004dffffffe6000000340000004e;
		5'b11011:	xpb = 256'h0000006c000000360000001b0000001b00000050ffffffe50000003600000051;
		5'b11100:	xpb = 256'h00000070000000380000001c0000001c00000053ffffffe40000003800000054;
		5'b11101:	xpb = 256'h000000740000003a0000001d0000001d00000056ffffffe30000003a00000057;
		5'b11110:	xpb = 256'h000000780000003c0000001e0000001e00000059ffffffe20000003c0000005a;
		5'b11111:	xpb = 256'h0000007c0000003e0000001f0000001f0000005cffffffe10000003e0000005d;
	endcase
end
endmodule

module xpb_32_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h000000800000004000000020000000200000005fffffffe00000004000000060;
		6'b000010:	xpb = 256'h00000100000000800000004000000040000000bfffffffc000000080000000c0;
		6'b000011:	xpb = 256'h00000180000000c000000060000000600000011fffffffa0000000c000000120;
		6'b000100:	xpb = 256'h000002000000010000000080000000800000017fffffff800000010000000180;
		6'b000101:	xpb = 256'h0000028000000140000000a0000000a0000001dfffffff6000000140000001e0;
		6'b000110:	xpb = 256'h0000030000000180000000c0000000c00000023fffffff400000018000000240;
		6'b000111:	xpb = 256'h00000380000001c0000000e0000000e00000029fffffff20000001c0000002a0;
		6'b001000:	xpb = 256'h00000400000002000000010000000100000002ffffffff000000020000000300;
		6'b001001:	xpb = 256'h000004800000024000000120000001200000035ffffffee00000024000000360;
		6'b001010:	xpb = 256'h00000500000002800000014000000140000003bffffffec000000280000003c0;
		6'b001011:	xpb = 256'h00000580000002c000000160000001600000041ffffffea0000002c000000420;
		6'b001100:	xpb = 256'h000006000000030000000180000001800000047ffffffe800000030000000480;
		6'b001101:	xpb = 256'h0000068000000340000001a0000001a0000004dffffffe6000000340000004e0;
		6'b001110:	xpb = 256'h0000070000000380000001c0000001c00000053ffffffe400000038000000540;
		6'b001111:	xpb = 256'h00000780000003c0000001e0000001e00000059ffffffe20000003c0000005a0;
		6'b010000:	xpb = 256'h00000800000004000000020000000200000005fffffffe000000040000000600;
		6'b010001:	xpb = 256'h000008800000044000000220000002200000065ffffffde00000044000000660;
		6'b010010:	xpb = 256'h00000900000004800000024000000240000006bffffffdc000000480000006c0;
		6'b010011:	xpb = 256'h00000980000004c000000260000002600000071ffffffda0000004c000000720;
		6'b010100:	xpb = 256'h00000a000000050000000280000002800000077ffffffd800000050000000780;
		6'b010101:	xpb = 256'h00000a8000000540000002a0000002a0000007dffffffd6000000540000007e0;
		6'b010110:	xpb = 256'h00000b0000000580000002c0000002c00000083ffffffd400000058000000840;
		6'b010111:	xpb = 256'h00000b80000005c0000002e0000002e00000089ffffffd20000005c0000008a0;
		6'b011000:	xpb = 256'h00000c00000006000000030000000300000008fffffffd000000060000000900;
		6'b011001:	xpb = 256'h00000c800000064000000320000003200000095ffffffce00000064000000960;
		6'b011010:	xpb = 256'h00000d00000006800000034000000340000009bffffffcc000000680000009c0;
		6'b011011:	xpb = 256'h00000d80000006c0000003600000036000000a1ffffffca0000006c000000a20;
		6'b011100:	xpb = 256'h00000e0000000700000003800000038000000a7ffffffc800000070000000a80;
		6'b011101:	xpb = 256'h00000e8000000740000003a0000003a000000adffffffc600000074000000ae0;
		6'b011110:	xpb = 256'h00000f0000000780000003c0000003c000000b3ffffffc400000078000000b40;
		6'b011111:	xpb = 256'h00000f80000007c0000003e0000003e000000b9ffffffc20000007c000000ba0;
		6'b100000:	xpb = 256'h0000100000000800000004000000040000000bfffffffc000000080000000c00;
		6'b100001:	xpb = 256'h0000108000000840000004200000042000000c5ffffffbe00000084000000c60;
		6'b100010:	xpb = 256'h0000110000000880000004400000044000000cbffffffbc00000088000000cc0;
		6'b100011:	xpb = 256'h00001180000008c0000004600000046000000d1ffffffba0000008c000000d20;
		6'b100100:	xpb = 256'h0000120000000900000004800000048000000d7ffffffb800000090000000d80;
		6'b100101:	xpb = 256'h0000128000000940000004a0000004a000000ddffffffb600000094000000de0;
		6'b100110:	xpb = 256'h0000130000000980000004c0000004c000000e3ffffffb400000098000000e40;
		6'b100111:	xpb = 256'h00001380000009c0000004e0000004e000000e9ffffffb20000009c000000ea0;
		6'b101000:	xpb = 256'h0000140000000a00000005000000050000000efffffffb0000000a0000000f00;
		6'b101001:	xpb = 256'h0000148000000a40000005200000052000000f5ffffffae000000a4000000f60;
		6'b101010:	xpb = 256'h0000150000000a80000005400000054000000fbffffffac000000a8000000fc0;
		6'b101011:	xpb = 256'h0000158000000ac000000560000005600000101ffffffaa000000ac000001020;
		6'b101100:	xpb = 256'h0000160000000b0000000580000005800000107ffffffa8000000b0000001080;
		6'b101101:	xpb = 256'h0000168000000b40000005a0000005a0000010dffffffa6000000b40000010e0;
		6'b101110:	xpb = 256'h0000170000000b80000005c0000005c00000113ffffffa4000000b8000001140;
		6'b101111:	xpb = 256'h0000178000000bc0000005e0000005e00000119ffffffa2000000bc0000011a0;
		6'b110000:	xpb = 256'h0000180000000c000000060000000600000011fffffffa0000000c0000001200;
		6'b110001:	xpb = 256'h0000188000000c4000000620000006200000125ffffff9e000000c4000001260;
		6'b110010:	xpb = 256'h0000190000000c800000064000000640000012bffffff9c000000c80000012c0;
		6'b110011:	xpb = 256'h0000198000000cc000000660000006600000131ffffff9a000000cc000001320;
		6'b110100:	xpb = 256'h00001a0000000d0000000680000006800000137ffffff98000000d0000001380;
		6'b110101:	xpb = 256'h00001a8000000d40000006a0000006a0000013dffffff96000000d40000013e0;
		6'b110110:	xpb = 256'h00001b0000000d80000006c0000006c00000143ffffff94000000d8000001440;
		6'b110111:	xpb = 256'h00001b8000000dc0000006e0000006e00000149ffffff92000000dc0000014a0;
		6'b111000:	xpb = 256'h00001c0000000e000000070000000700000014fffffff90000000e0000001500;
		6'b111001:	xpb = 256'h00001c8000000e4000000720000007200000155ffffff8e000000e4000001560;
		6'b111010:	xpb = 256'h00001d0000000e800000074000000740000015bffffff8c000000e80000015c0;
		6'b111011:	xpb = 256'h00001d8000000ec000000760000007600000161ffffff8a000000ec000001620;
		6'b111100:	xpb = 256'h00001e0000000f0000000780000007800000167ffffff88000000f0000001680;
		6'b111101:	xpb = 256'h00001e8000000f40000007a0000007a0000016dffffff86000000f40000016e0;
		6'b111110:	xpb = 256'h00001f0000000f80000007c0000007c00000173ffffff84000000f8000001740;
		6'b111111:	xpb = 256'h00001f8000000fc0000007e0000007e00000179ffffff82000000fc0000017a0;
	endcase
end
endmodule

module xpb_32_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00002000000010000000080000000800000017fffffff8000000100000001800;
		6'b000010:	xpb = 256'h0000400000002000000010000000100000002ffffffff0000000200000003000;
		6'b000011:	xpb = 256'h00006000000030000000180000001800000047ffffffe8000000300000004800;
		6'b000100:	xpb = 256'h0000800000004000000020000000200000005fffffffe0000000400000006000;
		6'b000101:	xpb = 256'h0000a000000050000000280000002800000077ffffffd8000000500000007800;
		6'b000110:	xpb = 256'h0000c00000006000000030000000300000008fffffffd0000000600000009000;
		6'b000111:	xpb = 256'h0000e0000000700000003800000038000000a7ffffffc800000070000000a800;
		6'b001000:	xpb = 256'h000100000000800000004000000040000000bfffffffc000000080000000c000;
		6'b001001:	xpb = 256'h000120000000900000004800000048000000d7ffffffb800000090000000d800;
		6'b001010:	xpb = 256'h000140000000a00000005000000050000000efffffffb0000000a0000000f000;
		6'b001011:	xpb = 256'h000160000000b0000000580000005800000107ffffffa8000000b00000010800;
		6'b001100:	xpb = 256'h000180000000c000000060000000600000011fffffffa0000000c00000012000;
		6'b001101:	xpb = 256'h0001a0000000d0000000680000006800000137ffffff98000000d00000013800;
		6'b001110:	xpb = 256'h0001c0000000e000000070000000700000014fffffff90000000e00000015000;
		6'b001111:	xpb = 256'h0001e0000000f0000000780000007800000167ffffff88000000f00000016800;
		6'b010000:	xpb = 256'h0002000000010000000080000000800000017fffffff80000001000000018000;
		6'b010001:	xpb = 256'h00022000000110000000880000008800000197ffffff78000001100000019800;
		6'b010010:	xpb = 256'h000240000001200000009000000090000001afffffff7000000120000001b000;
		6'b010011:	xpb = 256'h000260000001300000009800000098000001c7ffffff6800000130000001c800;
		6'b010100:	xpb = 256'h00028000000140000000a0000000a0000001dfffffff6000000140000001e000;
		6'b010101:	xpb = 256'h0002a000000150000000a8000000a8000001f7ffffff5800000150000001f800;
		6'b010110:	xpb = 256'h0002c000000160000000b0000000b00000020fffffff50000001600000021000;
		6'b010111:	xpb = 256'h0002e000000170000000b8000000b800000227ffffff48000001700000022800;
		6'b011000:	xpb = 256'h00030000000180000000c0000000c00000023fffffff40000001800000024000;
		6'b011001:	xpb = 256'h00032000000190000000c8000000c800000257ffffff38000001900000025800;
		6'b011010:	xpb = 256'h000340000001a0000000d0000000d00000026fffffff30000001a00000027000;
		6'b011011:	xpb = 256'h000360000001b0000000d8000000d800000287ffffff28000001b00000028800;
		6'b011100:	xpb = 256'h000380000001c0000000e0000000e00000029fffffff20000001c0000002a000;
		6'b011101:	xpb = 256'h0003a0000001d0000000e8000000e8000002b7ffffff18000001d0000002b800;
		6'b011110:	xpb = 256'h0003c0000001e0000000f0000000f0000002cfffffff10000001e0000002d000;
		6'b011111:	xpb = 256'h0003e0000001f0000000f8000000f8000002e7ffffff08000001f0000002e800;
		6'b100000:	xpb = 256'h000400000002000000010000000100000002ffffffff00000002000000030000;
		6'b100001:	xpb = 256'h00042000000210000001080000010800000317fffffef8000002100000031800;
		6'b100010:	xpb = 256'h0004400000022000000110000001100000032ffffffef0000002200000033000;
		6'b100011:	xpb = 256'h00046000000230000001180000011800000347fffffee8000002300000034800;
		6'b100100:	xpb = 256'h0004800000024000000120000001200000035ffffffee0000002400000036000;
		6'b100101:	xpb = 256'h0004a000000250000001280000012800000377fffffed8000002500000037800;
		6'b100110:	xpb = 256'h0004c00000026000000130000001300000038ffffffed0000002600000039000;
		6'b100111:	xpb = 256'h0004e0000002700000013800000138000003a7fffffec800000270000003a800;
		6'b101000:	xpb = 256'h000500000002800000014000000140000003bffffffec000000280000003c000;
		6'b101001:	xpb = 256'h000520000002900000014800000148000003d7fffffeb800000290000003d800;
		6'b101010:	xpb = 256'h000540000002a00000015000000150000003effffffeb0000002a0000003f000;
		6'b101011:	xpb = 256'h000560000002b0000001580000015800000407fffffea8000002b00000040800;
		6'b101100:	xpb = 256'h000580000002c000000160000001600000041ffffffea0000002c00000042000;
		6'b101101:	xpb = 256'h0005a0000002d0000001680000016800000437fffffe98000002d00000043800;
		6'b101110:	xpb = 256'h0005c0000002e000000170000001700000044ffffffe90000002e00000045000;
		6'b101111:	xpb = 256'h0005e0000002f0000001780000017800000467fffffe88000002f00000046800;
		6'b110000:	xpb = 256'h0006000000030000000180000001800000047ffffffe80000003000000048000;
		6'b110001:	xpb = 256'h00062000000310000001880000018800000497fffffe78000003100000049800;
		6'b110010:	xpb = 256'h000640000003200000019000000190000004affffffe7000000320000004b000;
		6'b110011:	xpb = 256'h000660000003300000019800000198000004c7fffffe6800000330000004c800;
		6'b110100:	xpb = 256'h00068000000340000001a0000001a0000004dffffffe6000000340000004e000;
		6'b110101:	xpb = 256'h0006a000000350000001a8000001a8000004f7fffffe5800000350000004f800;
		6'b110110:	xpb = 256'h0006c000000360000001b0000001b00000050ffffffe50000003600000051000;
		6'b110111:	xpb = 256'h0006e000000370000001b8000001b800000527fffffe48000003700000052800;
		6'b111000:	xpb = 256'h00070000000380000001c0000001c00000053ffffffe40000003800000054000;
		6'b111001:	xpb = 256'h00072000000390000001c8000001c800000557fffffe38000003900000055800;
		6'b111010:	xpb = 256'h000740000003a0000001d0000001d00000056ffffffe30000003a00000057000;
		6'b111011:	xpb = 256'h000760000003b0000001d8000001d800000587fffffe28000003b00000058800;
		6'b111100:	xpb = 256'h000780000003c0000001e0000001e00000059ffffffe20000003c0000005a000;
		6'b111101:	xpb = 256'h0007a0000003d0000001e8000001e8000005b7fffffe18000003d0000005b800;
		6'b111110:	xpb = 256'h0007c0000003e0000001f0000001f0000005cffffffe10000003e0000005d000;
		6'b111111:	xpb = 256'h0007e0000003f0000001f8000001f8000005e7fffffe08000003f0000005e800;
	endcase
end
endmodule

module xpb_33_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h000400000002000000010000000100000002ffffffff00000002000000030000;
		5'b00010:	xpb = 256'h000800000004000000020000000200000005fffffffe00000004000000060000;
		5'b00011:	xpb = 256'h000c00000006000000030000000300000008fffffffd00000006000000090000;
		5'b00100:	xpb = 256'h00100000000800000004000000040000000bfffffffc000000080000000c0000;
		5'b00101:	xpb = 256'h00140000000a00000005000000050000000efffffffb0000000a0000000f0000;
		5'b00110:	xpb = 256'h00180000000c000000060000000600000011fffffffa0000000c000000120000;
		5'b00111:	xpb = 256'h001c0000000e000000070000000700000014fffffff90000000e000000150000;
		5'b01000:	xpb = 256'h002000000010000000080000000800000017fffffff800000010000000180000;
		5'b01001:	xpb = 256'h00240000001200000009000000090000001afffffff7000000120000001b0000;
		5'b01010:	xpb = 256'h0028000000140000000a0000000a0000001dfffffff6000000140000001e0000;
		5'b01011:	xpb = 256'h002c000000160000000b0000000b00000020fffffff500000016000000210000;
		5'b01100:	xpb = 256'h0030000000180000000c0000000c00000023fffffff400000018000000240000;
		5'b01101:	xpb = 256'h00340000001a0000000d0000000d00000026fffffff30000001a000000270000;
		5'b01110:	xpb = 256'h00380000001c0000000e0000000e00000029fffffff20000001c0000002a0000;
		5'b01111:	xpb = 256'h003c0000001e0000000f0000000f0000002cfffffff10000001e0000002d0000;
		5'b10000:	xpb = 256'h00400000002000000010000000100000002ffffffff000000020000000300000;
		5'b10001:	xpb = 256'h004400000022000000110000001100000032ffffffef00000022000000330000;
		5'b10010:	xpb = 256'h004800000024000000120000001200000035ffffffee00000024000000360000;
		5'b10011:	xpb = 256'h004c00000026000000130000001300000038ffffffed00000026000000390000;
		5'b10100:	xpb = 256'h00500000002800000014000000140000003bffffffec000000280000003c0000;
		5'b10101:	xpb = 256'h00540000002a00000015000000150000003effffffeb0000002a0000003f0000;
		5'b10110:	xpb = 256'h00580000002c000000160000001600000041ffffffea0000002c000000420000;
		5'b10111:	xpb = 256'h005c0000002e000000170000001700000044ffffffe90000002e000000450000;
		5'b11000:	xpb = 256'h006000000030000000180000001800000047ffffffe800000030000000480000;
		5'b11001:	xpb = 256'h00640000003200000019000000190000004affffffe7000000320000004b0000;
		5'b11010:	xpb = 256'h0068000000340000001a0000001a0000004dffffffe6000000340000004e0000;
		5'b11011:	xpb = 256'h006c000000360000001b0000001b00000050ffffffe500000036000000510000;
		5'b11100:	xpb = 256'h0070000000380000001c0000001c00000053ffffffe400000038000000540000;
		5'b11101:	xpb = 256'h00740000003a0000001d0000001d00000056ffffffe30000003a000000570000;
		5'b11110:	xpb = 256'h00780000003c0000001e0000001e00000059ffffffe20000003c0000005a0000;
		5'b11111:	xpb = 256'h007c0000003e0000001f0000001f0000005cffffffe10000003e0000005d0000;
	endcase
end
endmodule

module xpb_33_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00800000004000000020000000200000005fffffffe000000040000000600000;
		6'b000010:	xpb = 256'h0100000000800000004000000040000000bfffffffc000000080000000c00000;
		6'b000011:	xpb = 256'h0180000000c000000060000000600000011fffffffa0000000c0000001200000;
		6'b000100:	xpb = 256'h02000000010000000080000000800000017fffffff8000000100000001800000;
		6'b000101:	xpb = 256'h028000000140000000a0000000a0000001dfffffff6000000140000001e00000;
		6'b000110:	xpb = 256'h030000000180000000c0000000c00000023fffffff4000000180000002400000;
		6'b000111:	xpb = 256'h0380000001c0000000e0000000e00000029fffffff20000001c0000002a00000;
		6'b001000:	xpb = 256'h0400000002000000010000000100000002ffffffff0000000200000003000000;
		6'b001001:	xpb = 256'h04800000024000000120000001200000035ffffffee000000240000003600000;
		6'b001010:	xpb = 256'h0500000002800000014000000140000003bffffffec000000280000003c00000;
		6'b001011:	xpb = 256'h0580000002c000000160000001600000041ffffffea0000002c0000004200000;
		6'b001100:	xpb = 256'h06000000030000000180000001800000047ffffffe8000000300000004800000;
		6'b001101:	xpb = 256'h068000000340000001a0000001a0000004dffffffe6000000340000004e00000;
		6'b001110:	xpb = 256'h070000000380000001c0000001c00000053ffffffe4000000380000005400000;
		6'b001111:	xpb = 256'h0780000003c0000001e0000001e00000059ffffffe20000003c0000005a00000;
		6'b010000:	xpb = 256'h0800000004000000020000000200000005fffffffe0000000400000006000000;
		6'b010001:	xpb = 256'h08800000044000000220000002200000065ffffffde000000440000006600000;
		6'b010010:	xpb = 256'h0900000004800000024000000240000006bffffffdc000000480000006c00000;
		6'b010011:	xpb = 256'h0980000004c000000260000002600000071ffffffda0000004c0000007200000;
		6'b010100:	xpb = 256'h0a000000050000000280000002800000077ffffffd8000000500000007800000;
		6'b010101:	xpb = 256'h0a8000000540000002a0000002a0000007dffffffd6000000540000007e00000;
		6'b010110:	xpb = 256'h0b0000000580000002c0000002c00000083ffffffd4000000580000008400000;
		6'b010111:	xpb = 256'h0b80000005c0000002e0000002e00000089ffffffd20000005c0000008a00000;
		6'b011000:	xpb = 256'h0c00000006000000030000000300000008fffffffd0000000600000009000000;
		6'b011001:	xpb = 256'h0c800000064000000320000003200000095ffffffce000000640000009600000;
		6'b011010:	xpb = 256'h0d00000006800000034000000340000009bffffffcc000000680000009c00000;
		6'b011011:	xpb = 256'h0d80000006c0000003600000036000000a1ffffffca0000006c000000a200000;
		6'b011100:	xpb = 256'h0e0000000700000003800000038000000a7ffffffc800000070000000a800000;
		6'b011101:	xpb = 256'h0e8000000740000003a0000003a000000adffffffc600000074000000ae00000;
		6'b011110:	xpb = 256'h0f0000000780000003c0000003c000000b3ffffffc400000078000000b400000;
		6'b011111:	xpb = 256'h0f80000007c0000003e0000003e000000b9ffffffc20000007c000000ba00000;
		6'b100000:	xpb = 256'h100000000800000004000000040000000bfffffffc000000080000000c000000;
		6'b100001:	xpb = 256'h108000000840000004200000042000000c5ffffffbe00000084000000c600000;
		6'b100010:	xpb = 256'h110000000880000004400000044000000cbffffffbc00000088000000cc00000;
		6'b100011:	xpb = 256'h1180000008c0000004600000046000000d1ffffffba0000008c000000d200000;
		6'b100100:	xpb = 256'h120000000900000004800000048000000d7ffffffb800000090000000d800000;
		6'b100101:	xpb = 256'h128000000940000004a0000004a000000ddffffffb600000094000000de00000;
		6'b100110:	xpb = 256'h130000000980000004c0000004c000000e3ffffffb400000098000000e400000;
		6'b100111:	xpb = 256'h1380000009c0000004e0000004e000000e9ffffffb20000009c000000ea00000;
		6'b101000:	xpb = 256'h140000000a00000005000000050000000efffffffb0000000a0000000f000000;
		6'b101001:	xpb = 256'h148000000a40000005200000052000000f5ffffffae000000a4000000f600000;
		6'b101010:	xpb = 256'h150000000a80000005400000054000000fbffffffac000000a8000000fc00000;
		6'b101011:	xpb = 256'h158000000ac000000560000005600000101ffffffaa000000ac0000010200000;
		6'b101100:	xpb = 256'h160000000b0000000580000005800000107ffffffa8000000b00000010800000;
		6'b101101:	xpb = 256'h168000000b40000005a0000005a0000010dffffffa6000000b40000010e00000;
		6'b101110:	xpb = 256'h170000000b80000005c0000005c00000113ffffffa4000000b80000011400000;
		6'b101111:	xpb = 256'h178000000bc0000005e0000005e00000119ffffffa2000000bc0000011a00000;
		6'b110000:	xpb = 256'h180000000c000000060000000600000011fffffffa0000000c00000012000000;
		6'b110001:	xpb = 256'h188000000c4000000620000006200000125ffffff9e000000c40000012600000;
		6'b110010:	xpb = 256'h190000000c800000064000000640000012bffffff9c000000c80000012c00000;
		6'b110011:	xpb = 256'h198000000cc000000660000006600000131ffffff9a000000cc0000013200000;
		6'b110100:	xpb = 256'h1a0000000d0000000680000006800000137ffffff98000000d00000013800000;
		6'b110101:	xpb = 256'h1a8000000d40000006a0000006a0000013dffffff96000000d40000013e00000;
		6'b110110:	xpb = 256'h1b0000000d80000006c0000006c00000143ffffff94000000d80000014400000;
		6'b110111:	xpb = 256'h1b8000000dc0000006e0000006e00000149ffffff92000000dc0000014a00000;
		6'b111000:	xpb = 256'h1c0000000e000000070000000700000014fffffff90000000e00000015000000;
		6'b111001:	xpb = 256'h1c8000000e4000000720000007200000155ffffff8e000000e40000015600000;
		6'b111010:	xpb = 256'h1d0000000e800000074000000740000015bffffff8c000000e80000015c00000;
		6'b111011:	xpb = 256'h1d8000000ec000000760000007600000161ffffff8a000000ec0000016200000;
		6'b111100:	xpb = 256'h1e0000000f0000000780000007800000167ffffff88000000f00000016800000;
		6'b111101:	xpb = 256'h1e8000000f40000007a0000007a0000016dffffff86000000f40000016e00000;
		6'b111110:	xpb = 256'h1f0000000f80000007c0000007c00000173ffffff84000000f80000017400000;
		6'b111111:	xpb = 256'h1f8000000fc0000007e0000007e00000179ffffff82000000fc0000017a00000;
	endcase
end
endmodule

module xpb_33_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h2000000010000000080000000800000017fffffff80000001000000018000000;
		6'b000010:	xpb = 256'h400000002000000010000000100000002ffffffff00000002000000030000000;
		6'b000011:	xpb = 256'h6000000030000000180000001800000047ffffffe80000003000000048000000;
		6'b000100:	xpb = 256'h800000004000000020000000200000005fffffffe00000004000000060000000;
		6'b000101:	xpb = 256'ha000000050000000280000002800000077ffffffd80000005000000078000000;
		6'b000110:	xpb = 256'hc00000006000000030000000300000008fffffffd00000006000000090000000;
		6'b000111:	xpb = 256'he0000000700000003800000038000000a7ffffffc800000070000000a8000000;
		6'b001000:	xpb = 256'h00000001800000004000000040000000c0000000bfffffff80000000c0000001;
		6'b001001:	xpb = 256'h20000001900000004800000048000000d8000000b7ffffff90000000d8000001;
		6'b001010:	xpb = 256'h40000001a00000005000000050000000f0000000afffffffa0000000f0000001;
		6'b001011:	xpb = 256'h60000001b0000000580000005800000108000000a7ffffffb000000108000001;
		6'b001100:	xpb = 256'h80000001c00000006000000060000001200000009fffffffc000000120000001;
		6'b001101:	xpb = 256'ha0000001d000000068000000680000013800000097ffffffd000000138000001;
		6'b001110:	xpb = 256'hc0000001e00000007000000070000001500000008fffffffe000000150000001;
		6'b001111:	xpb = 256'he0000001f000000078000000780000016800000087fffffff000000168000001;
		6'b010000:	xpb = 256'h00000003000000008000000080000001800000017fffffff0000000180000002;
		6'b010001:	xpb = 256'h200000031000000088000000880000019800000177ffffff1000000198000002;
		6'b010010:	xpb = 256'h40000003200000009000000090000001b00000016fffffff20000001b0000002;
		6'b010011:	xpb = 256'h60000003300000009800000098000001c800000167ffffff30000001c8000002;
		6'b010100:	xpb = 256'h8000000340000000a0000000a0000001e00000015fffffff40000001e0000002;
		6'b010101:	xpb = 256'ha000000350000000a8000000a8000001f800000157ffffff50000001f8000002;
		6'b010110:	xpb = 256'hc000000360000000b0000000b0000002100000014fffffff6000000210000002;
		6'b010111:	xpb = 256'he000000370000000b8000000b80000022800000147ffffff7000000228000002;
		6'b011000:	xpb = 256'h0000000480000000c0000000c0000002400000023ffffffe8000000240000003;
		6'b011001:	xpb = 256'h2000000490000000c8000000c80000025800000237fffffe9000000258000003;
		6'b011010:	xpb = 256'h40000004a0000000d0000000d0000002700000022ffffffea000000270000003;
		6'b011011:	xpb = 256'h60000004b0000000d8000000d80000028800000227fffffeb000000288000003;
		6'b011100:	xpb = 256'h80000004c0000000e0000000e0000002a00000021ffffffec0000002a0000003;
		6'b011101:	xpb = 256'ha0000004d0000000e8000000e8000002b800000217fffffed0000002b8000003;
		6'b011110:	xpb = 256'hc0000004e0000000f0000000f0000002d00000020ffffffee0000002d0000003;
		6'b011111:	xpb = 256'he0000004f0000000f8000000f8000002e800000207fffffef0000002e8000003;
		6'b100000:	xpb = 256'h0000000600000001000000010000000300000002fffffffe0000000300000004;
		6'b100001:	xpb = 256'h2000000610000001080000010800000318000002f7fffffe1000000318000004;
		6'b100010:	xpb = 256'h4000000620000001100000011000000330000002effffffe2000000330000004;
		6'b100011:	xpb = 256'h6000000630000001180000011800000348000002e7fffffe3000000348000004;
		6'b100100:	xpb = 256'h8000000640000001200000012000000360000002dffffffe4000000360000004;
		6'b100101:	xpb = 256'ha000000650000001280000012800000378000002d7fffffe5000000378000004;
		6'b100110:	xpb = 256'hc000000660000001300000013000000390000002cffffffe6000000390000004;
		6'b100111:	xpb = 256'he0000006700000013800000138000003a8000002c7fffffe70000003a8000004;
		6'b101000:	xpb = 256'h00000007800000014000000140000003c0000003bffffffd80000003c0000005;
		6'b101001:	xpb = 256'h20000007900000014800000148000003d8000003b7fffffd90000003d8000005;
		6'b101010:	xpb = 256'h40000007a00000015000000150000003f0000003affffffda0000003f0000005;
		6'b101011:	xpb = 256'h60000007b0000001580000015800000408000003a7fffffdb000000408000005;
		6'b101100:	xpb = 256'h80000007c00000016000000160000004200000039ffffffdc000000420000005;
		6'b101101:	xpb = 256'ha0000007d000000168000001680000043800000397fffffdd000000438000005;
		6'b101110:	xpb = 256'hc0000007e00000017000000170000004500000038ffffffde000000450000005;
		6'b101111:	xpb = 256'he0000007f000000178000001780000046800000387fffffdf000000468000005;
		6'b110000:	xpb = 256'h00000009000000018000000180000004800000047ffffffd0000000480000006;
		6'b110001:	xpb = 256'h200000091000000188000001880000049800000477fffffd1000000498000006;
		6'b110010:	xpb = 256'h40000009200000019000000190000004b00000046ffffffd20000004b0000006;
		6'b110011:	xpb = 256'h60000009300000019800000198000004c800000467fffffd30000004c8000006;
		6'b110100:	xpb = 256'h8000000940000001a0000001a0000004e00000045ffffffd40000004e0000006;
		6'b110101:	xpb = 256'ha000000950000001a8000001a8000004f800000457fffffd50000004f8000006;
		6'b110110:	xpb = 256'hc000000960000001b0000001b0000005100000044ffffffd6000000510000006;
		6'b110111:	xpb = 256'he000000970000001b8000001b80000052800000447fffffd7000000528000006;
		6'b111000:	xpb = 256'h0000000a80000001c0000001c0000005400000053ffffffc8000000540000007;
		6'b111001:	xpb = 256'h2000000a90000001c8000001c80000055800000537fffffc9000000558000007;
		6'b111010:	xpb = 256'h4000000aa0000001d0000001d0000005700000052ffffffca000000570000007;
		6'b111011:	xpb = 256'h6000000ab0000001d8000001d80000058800000527fffffcb000000588000007;
		6'b111100:	xpb = 256'h8000000ac0000001e0000001e0000005a00000051ffffffcc0000005a0000007;
		6'b111101:	xpb = 256'ha000000ad0000001e8000001e8000005b800000517fffffcd0000005b8000007;
		6'b111110:	xpb = 256'hc000000ae0000001f0000001f0000005d00000050ffffffce0000005d0000007;
		6'b111111:	xpb = 256'he000000af0000001f8000001f8000005e800000507fffffcf0000005e8000007;
	endcase
end
endmodule

module xpb_34_lsb
(
    input logic [4:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		5'b00000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		5'b00001:	xpb = 256'h0000000600000001000000010000000300000002fffffffe0000000300000004;
		5'b00010:	xpb = 256'h0000000c00000002000000020000000600000005fffffffc0000000600000008;
		5'b00011:	xpb = 256'h0000001200000003000000030000000900000008fffffffa000000090000000c;
		5'b00100:	xpb = 256'h0000001800000004000000040000000c0000000bfffffff80000000c00000010;
		5'b00101:	xpb = 256'h0000001e00000005000000050000000f0000000efffffff60000000f00000014;
		5'b00110:	xpb = 256'h0000002400000006000000060000001200000011fffffff40000001200000018;
		5'b00111:	xpb = 256'h0000002a00000007000000070000001500000014fffffff2000000150000001c;
		5'b01000:	xpb = 256'h0000003000000008000000080000001800000017fffffff00000001800000020;
		5'b01001:	xpb = 256'h0000003600000009000000090000001b0000001affffffee0000001b00000024;
		5'b01010:	xpb = 256'h0000003c0000000a0000000a0000001e0000001dffffffec0000001e00000028;
		5'b01011:	xpb = 256'h000000420000000b0000000b0000002100000020ffffffea000000210000002c;
		5'b01100:	xpb = 256'h000000480000000c0000000c0000002400000023ffffffe80000002400000030;
		5'b01101:	xpb = 256'h0000004e0000000d0000000d0000002700000026ffffffe60000002700000034;
		5'b01110:	xpb = 256'h000000540000000e0000000e0000002a00000029ffffffe40000002a00000038;
		5'b01111:	xpb = 256'h0000005a0000000f0000000f0000002d0000002cffffffe20000002d0000003c;
		5'b10000:	xpb = 256'h000000600000001000000010000000300000002fffffffe00000003000000040;
		5'b10001:	xpb = 256'h0000006600000011000000110000003300000032ffffffde0000003300000044;
		5'b10010:	xpb = 256'h0000006c00000012000000120000003600000035ffffffdc0000003600000048;
		5'b10011:	xpb = 256'h0000007200000013000000130000003900000038ffffffda000000390000004c;
		5'b10100:	xpb = 256'h0000007800000014000000140000003c0000003bffffffd80000003c00000050;
		5'b10101:	xpb = 256'h0000007e00000015000000150000003f0000003effffffd60000003f00000054;
		5'b10110:	xpb = 256'h0000008400000016000000160000004200000041ffffffd40000004200000058;
		5'b10111:	xpb = 256'h0000008a00000017000000170000004500000044ffffffd2000000450000005c;
		5'b11000:	xpb = 256'h0000009000000018000000180000004800000047ffffffd00000004800000060;
		5'b11001:	xpb = 256'h0000009600000019000000190000004b0000004affffffce0000004b00000064;
		5'b11010:	xpb = 256'h0000009c0000001a0000001a0000004e0000004dffffffcc0000004e00000068;
		5'b11011:	xpb = 256'h000000a20000001b0000001b0000005100000050ffffffca000000510000006c;
		5'b11100:	xpb = 256'h000000a80000001c0000001c0000005400000053ffffffc80000005400000070;
		5'b11101:	xpb = 256'h000000ae0000001d0000001d0000005700000056ffffffc60000005700000074;
		5'b11110:	xpb = 256'h000000b40000001e0000001e0000005a00000059ffffffc40000005a00000078;
		5'b11111:	xpb = 256'h000000ba0000001f0000001f0000005d0000005cffffffc20000005d0000007c;
	endcase
end
endmodule

module xpb_34_csb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h000000c00000002000000020000000600000005fffffffc00000006000000080;
		6'b000010:	xpb = 256'h000001800000004000000040000000c0000000bfffffff80000000c000000100;
		6'b000011:	xpb = 256'h000002400000006000000060000001200000011fffffff400000012000000180;
		6'b000100:	xpb = 256'h000003000000008000000080000001800000017fffffff000000018000000200;
		6'b000101:	xpb = 256'h000003c0000000a0000000a0000001e0000001dffffffec0000001e000000280;
		6'b000110:	xpb = 256'h00000480000000c0000000c0000002400000023ffffffe800000024000000300;
		6'b000111:	xpb = 256'h00000540000000e0000000e0000002a00000029ffffffe40000002a000000380;
		6'b001000:	xpb = 256'h00000600000001000000010000000300000002fffffffe000000030000000400;
		6'b001001:	xpb = 256'h000006c00000012000000120000003600000035ffffffdc00000036000000480;
		6'b001010:	xpb = 256'h000007800000014000000140000003c0000003bffffffd80000003c000000500;
		6'b001011:	xpb = 256'h000008400000016000000160000004200000041ffffffd400000042000000580;
		6'b001100:	xpb = 256'h000009000000018000000180000004800000047ffffffd000000048000000600;
		6'b001101:	xpb = 256'h000009c0000001a0000001a0000004e0000004dffffffcc0000004e000000680;
		6'b001110:	xpb = 256'h00000a80000001c0000001c0000005400000053ffffffc800000054000000700;
		6'b001111:	xpb = 256'h00000b40000001e0000001e0000005a00000059ffffffc40000005a000000780;
		6'b010000:	xpb = 256'h00000c00000002000000020000000600000005fffffffc000000060000000800;
		6'b010001:	xpb = 256'h00000cc00000022000000220000006600000065ffffffbc00000066000000880;
		6'b010010:	xpb = 256'h00000d800000024000000240000006c0000006bffffffb80000006c000000900;
		6'b010011:	xpb = 256'h00000e400000026000000260000007200000071ffffffb400000072000000980;
		6'b010100:	xpb = 256'h00000f000000028000000280000007800000077ffffffb000000078000000a00;
		6'b010101:	xpb = 256'h00000fc0000002a0000002a0000007e0000007dffffffac0000007e000000a80;
		6'b010110:	xpb = 256'h00001080000002c0000002c0000008400000083ffffffa800000084000000b00;
		6'b010111:	xpb = 256'h00001140000002e0000002e0000008a00000089ffffffa40000008a000000b80;
		6'b011000:	xpb = 256'h00001200000003000000030000000900000008fffffffa000000090000000c00;
		6'b011001:	xpb = 256'h000012c00000032000000320000009600000095ffffff9c00000096000000c80;
		6'b011010:	xpb = 256'h000013800000034000000340000009c0000009bffffff980000009c000000d00;
		6'b011011:	xpb = 256'h00001440000003600000036000000a2000000a1ffffff94000000a2000000d80;
		6'b011100:	xpb = 256'h00001500000003800000038000000a8000000a7ffffff90000000a8000000e00;
		6'b011101:	xpb = 256'h000015c0000003a0000003a000000ae000000adffffff8c000000ae000000e80;
		6'b011110:	xpb = 256'h00001680000003c0000003c000000b4000000b3ffffff88000000b4000000f00;
		6'b011111:	xpb = 256'h00001740000003e0000003e000000ba000000b9ffffff84000000ba000000f80;
		6'b100000:	xpb = 256'h00001800000004000000040000000c0000000bfffffff80000000c0000001000;
		6'b100001:	xpb = 256'h000018c0000004200000042000000c6000000c5ffffff7c000000c6000001080;
		6'b100010:	xpb = 256'h00001980000004400000044000000cc000000cbffffff78000000cc000001100;
		6'b100011:	xpb = 256'h00001a40000004600000046000000d2000000d1ffffff74000000d2000001180;
		6'b100100:	xpb = 256'h00001b00000004800000048000000d8000000d7ffffff70000000d8000001200;
		6'b100101:	xpb = 256'h00001bc0000004a0000004a000000de000000ddffffff6c000000de000001280;
		6'b100110:	xpb = 256'h00001c80000004c0000004c000000e4000000e3ffffff68000000e4000001300;
		6'b100111:	xpb = 256'h00001d40000004e0000004e000000ea000000e9ffffff64000000ea000001380;
		6'b101000:	xpb = 256'h00001e00000005000000050000000f0000000efffffff60000000f0000001400;
		6'b101001:	xpb = 256'h00001ec0000005200000052000000f6000000f5ffffff5c000000f6000001480;
		6'b101010:	xpb = 256'h00001f80000005400000054000000fc000000fbffffff58000000fc000001500;
		6'b101011:	xpb = 256'h000020400000056000000560000010200000101ffffff5400000102000001580;
		6'b101100:	xpb = 256'h000021000000058000000580000010800000107ffffff5000000108000001600;
		6'b101101:	xpb = 256'h000021c0000005a0000005a0000010e0000010dffffff4c0000010e000001680;
		6'b101110:	xpb = 256'h00002280000005c0000005c0000011400000113ffffff4800000114000001700;
		6'b101111:	xpb = 256'h00002340000005e0000005e0000011a00000119ffffff440000011a000001780;
		6'b110000:	xpb = 256'h00002400000006000000060000001200000011fffffff4000000120000001800;
		6'b110001:	xpb = 256'h000024c00000062000000620000012600000125ffffff3c00000126000001880;
		6'b110010:	xpb = 256'h000025800000064000000640000012c0000012bffffff380000012c000001900;
		6'b110011:	xpb = 256'h000026400000066000000660000013200000131ffffff3400000132000001980;
		6'b110100:	xpb = 256'h000027000000068000000680000013800000137ffffff3000000138000001a00;
		6'b110101:	xpb = 256'h000027c0000006a0000006a0000013e0000013dffffff2c0000013e000001a80;
		6'b110110:	xpb = 256'h00002880000006c0000006c0000014400000143ffffff2800000144000001b00;
		6'b110111:	xpb = 256'h00002940000006e0000006e0000014a00000149ffffff240000014a000001b80;
		6'b111000:	xpb = 256'h00002a00000007000000070000001500000014fffffff2000000150000001c00;
		6'b111001:	xpb = 256'h00002ac00000072000000720000015600000155ffffff1c00000156000001c80;
		6'b111010:	xpb = 256'h00002b800000074000000740000015c0000015bffffff180000015c000001d00;
		6'b111011:	xpb = 256'h00002c400000076000000760000016200000161ffffff1400000162000001d80;
		6'b111100:	xpb = 256'h00002d000000078000000780000016800000167ffffff1000000168000001e00;
		6'b111101:	xpb = 256'h00002dc0000007a0000007a0000016e0000016dffffff0c0000016e000001e80;
		6'b111110:	xpb = 256'h00002e80000007c0000007c0000017400000173ffffff0800000174000001f00;
		6'b111111:	xpb = 256'h00002f40000007e0000007e0000017a00000179ffffff040000017a000001f80;
	endcase
end
endmodule

module xpb_34_msb
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h00003000000008000000080000001800000017fffffff0000000180000002000;
		6'b000010:	xpb = 256'h0000600000001000000010000000300000002fffffffe0000000300000004000;
		6'b000011:	xpb = 256'h00009000000018000000180000004800000047ffffffd0000000480000006000;
		6'b000100:	xpb = 256'h0000c00000002000000020000000600000005fffffffc0000000600000008000;
		6'b000101:	xpb = 256'h0000f000000028000000280000007800000077ffffffb000000078000000a000;
		6'b000110:	xpb = 256'h0001200000003000000030000000900000008fffffffa000000090000000c000;
		6'b000111:	xpb = 256'h0001500000003800000038000000a8000000a7ffffff90000000a8000000e000;
		6'b001000:	xpb = 256'h0001800000004000000040000000c0000000bfffffff80000000c00000010000;
		6'b001001:	xpb = 256'h0001b00000004800000048000000d8000000d7ffffff70000000d80000012000;
		6'b001010:	xpb = 256'h0001e00000005000000050000000f0000000efffffff60000000f00000014000;
		6'b001011:	xpb = 256'h00021000000058000000580000010800000107ffffff50000001080000016000;
		6'b001100:	xpb = 256'h0002400000006000000060000001200000011fffffff40000001200000018000;
		6'b001101:	xpb = 256'h00027000000068000000680000013800000137ffffff3000000138000001a000;
		6'b001110:	xpb = 256'h0002a00000007000000070000001500000014fffffff2000000150000001c000;
		6'b001111:	xpb = 256'h0002d000000078000000780000016800000167ffffff1000000168000001e000;
		6'b010000:	xpb = 256'h0003000000008000000080000001800000017fffffff00000001800000020000;
		6'b010001:	xpb = 256'h00033000000088000000880000019800000197fffffef0000001980000022000;
		6'b010010:	xpb = 256'h0003600000009000000090000001b0000001affffffee0000001b00000024000;
		6'b010011:	xpb = 256'h0003900000009800000098000001c8000001c7fffffed0000001c80000026000;
		6'b010100:	xpb = 256'h0003c0000000a0000000a0000001e0000001dffffffec0000001e00000028000;
		6'b010101:	xpb = 256'h0003f0000000a8000000a8000001f8000001f7fffffeb0000001f8000002a000;
		6'b010110:	xpb = 256'h000420000000b0000000b0000002100000020ffffffea000000210000002c000;
		6'b010111:	xpb = 256'h000450000000b8000000b80000022800000227fffffe9000000228000002e000;
		6'b011000:	xpb = 256'h000480000000c0000000c0000002400000023ffffffe80000002400000030000;
		6'b011001:	xpb = 256'h0004b0000000c8000000c80000025800000257fffffe70000002580000032000;
		6'b011010:	xpb = 256'h0004e0000000d0000000d0000002700000026ffffffe60000002700000034000;
		6'b011011:	xpb = 256'h000510000000d8000000d80000028800000287fffffe50000002880000036000;
		6'b011100:	xpb = 256'h000540000000e0000000e0000002a00000029ffffffe40000002a00000038000;
		6'b011101:	xpb = 256'h000570000000e8000000e8000002b8000002b7fffffe30000002b8000003a000;
		6'b011110:	xpb = 256'h0005a0000000f0000000f0000002d0000002cffffffe20000002d0000003c000;
		6'b011111:	xpb = 256'h0005d0000000f8000000f8000002e8000002e7fffffe10000002e8000003e000;
		6'b100000:	xpb = 256'h000600000001000000010000000300000002fffffffe00000003000000040000;
		6'b100001:	xpb = 256'h00063000000108000001080000031800000317fffffdf0000003180000042000;
		6'b100010:	xpb = 256'h0006600000011000000110000003300000032ffffffde0000003300000044000;
		6'b100011:	xpb = 256'h00069000000118000001180000034800000347fffffdd0000003480000046000;
		6'b100100:	xpb = 256'h0006c00000012000000120000003600000035ffffffdc0000003600000048000;
		6'b100101:	xpb = 256'h0006f000000128000001280000037800000377fffffdb000000378000004a000;
		6'b100110:	xpb = 256'h0007200000013000000130000003900000038ffffffda000000390000004c000;
		6'b100111:	xpb = 256'h0007500000013800000138000003a8000003a7fffffd90000003a8000004e000;
		6'b101000:	xpb = 256'h0007800000014000000140000003c0000003bffffffd80000003c00000050000;
		6'b101001:	xpb = 256'h0007b00000014800000148000003d8000003d7fffffd70000003d80000052000;
		6'b101010:	xpb = 256'h0007e00000015000000150000003f0000003effffffd60000003f00000054000;
		6'b101011:	xpb = 256'h00081000000158000001580000040800000407fffffd50000004080000056000;
		6'b101100:	xpb = 256'h0008400000016000000160000004200000041ffffffd40000004200000058000;
		6'b101101:	xpb = 256'h00087000000168000001680000043800000437fffffd3000000438000005a000;
		6'b101110:	xpb = 256'h0008a00000017000000170000004500000044ffffffd2000000450000005c000;
		6'b101111:	xpb = 256'h0008d000000178000001780000046800000467fffffd1000000468000005e000;
		6'b110000:	xpb = 256'h0009000000018000000180000004800000047ffffffd00000004800000060000;
		6'b110001:	xpb = 256'h00093000000188000001880000049800000497fffffcf0000004980000062000;
		6'b110010:	xpb = 256'h0009600000019000000190000004b0000004affffffce0000004b00000064000;
		6'b110011:	xpb = 256'h0009900000019800000198000004c8000004c7fffffcd0000004c80000066000;
		6'b110100:	xpb = 256'h0009c0000001a0000001a0000004e0000004dffffffcc0000004e00000068000;
		6'b110101:	xpb = 256'h0009f0000001a8000001a8000004f8000004f7fffffcb0000004f8000006a000;
		6'b110110:	xpb = 256'h000a20000001b0000001b0000005100000050ffffffca000000510000006c000;
		6'b110111:	xpb = 256'h000a50000001b8000001b80000052800000527fffffc9000000528000006e000;
		6'b111000:	xpb = 256'h000a80000001c0000001c0000005400000053ffffffc80000005400000070000;
		6'b111001:	xpb = 256'h000ab0000001c8000001c80000055800000557fffffc70000005580000072000;
		6'b111010:	xpb = 256'h000ae0000001d0000001d0000005700000056ffffffc60000005700000074000;
		6'b111011:	xpb = 256'h000b10000001d8000001d80000058800000587fffffc50000005880000076000;
		6'b111100:	xpb = 256'h000b40000001e0000001e0000005a00000059ffffffc40000005a00000078000;
		6'b111101:	xpb = 256'h000b70000001e8000001e8000005b8000005b7fffffc30000005b8000007a000;
		6'b111110:	xpb = 256'h000ba0000001f0000001f0000005d0000005cffffffc20000005d0000007c000;
		6'b111111:	xpb = 256'h000bd0000001f8000001f8000005e8000005e7fffffc10000005e8000007e000;
	endcase
end
endmodule
