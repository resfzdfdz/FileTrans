/*******************************************************************************
  Copyright 2019 Xi'an Jiaotong University

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
*******************************************************************************/

module xpb_addsub
(
    input logic [5:0]          x,
    output logic [15:0] [15:0] xpb
);

always_comb begin
    case(x)
		6'b000000:	xpb = 256'h0000000000000000000000000000000000000000000000000000000000000000;
		6'b000001:	xpb = 256'h0000000100000000000000000000000000000000ffffffff0000000000000001;
		6'b000010:	xpb = 256'h0000000200000000000000000000000000000001fffffffe0000000000000002;
		6'b000011:	xpb = 256'h0000000300000000000000000000000000000002fffffffd0000000000000003;
		6'b000100:	xpb = 256'h0000000400000000000000000000000000000003fffffffc0000000000000004;
		6'b000101:	xpb = 256'h0000000500000000000000000000000000000004fffffffb0000000000000005;
		6'b000110:	xpb = 256'h0000000600000000000000000000000000000005fffffffa0000000000000006;
		6'b000111:	xpb = 256'h0000000700000000000000000000000000000006fffffff90000000000000007;
		6'b001000:	xpb = 256'h0000000800000000000000000000000000000007fffffff80000000000000008;
		6'b001001:	xpb = 256'h0000000900000000000000000000000000000008fffffff70000000000000009;
		6'b001010:	xpb = 256'h0000000a00000000000000000000000000000009fffffff6000000000000000a;
		6'b001011:	xpb = 256'h0000000b0000000000000000000000000000000afffffff5000000000000000b;
		6'b001100:	xpb = 256'h0000000c0000000000000000000000000000000bfffffff4000000000000000c;
		6'b001101:	xpb = 256'h0000000d0000000000000000000000000000000cfffffff3000000000000000d;
		6'b001110:	xpb = 256'h0000000e0000000000000000000000000000000dfffffff2000000000000000e;
		6'b001111:	xpb = 256'h0000000f0000000000000000000000000000000efffffff1000000000000000f;
		6'b010000:	xpb = 256'h000000100000000000000000000000000000000ffffffff00000000000000010;
		6'b010001:	xpb = 256'h0000001100000000000000000000000000000010ffffffef0000000000000011;
		6'b010010:	xpb = 256'h0000001200000000000000000000000000000011ffffffee0000000000000012;
		6'b010011:	xpb = 256'h0000001300000000000000000000000000000012ffffffed0000000000000013;
		6'b010100:	xpb = 256'h0000001400000000000000000000000000000013ffffffec0000000000000014;
		6'b010101:	xpb = 256'h0000001500000000000000000000000000000014ffffffeb0000000000000015;
		6'b010110:	xpb = 256'h0000001600000000000000000000000000000015ffffffea0000000000000016;
		6'b010111:	xpb = 256'h0000001700000000000000000000000000000016ffffffe90000000000000017;
		6'b011000:	xpb = 256'h0000001800000000000000000000000000000017ffffffe80000000000000018;
		6'b011001:	xpb = 256'h0000001900000000000000000000000000000018ffffffe70000000000000019;
		6'b011010:	xpb = 256'h0000001a00000000000000000000000000000019ffffffe6000000000000001a;
		6'b011011:	xpb = 256'h0000001b0000000000000000000000000000001affffffe5000000000000001b;
		6'b011100:	xpb = 256'h0000001c0000000000000000000000000000001bffffffe4000000000000001c;
		6'b011101:	xpb = 256'h0000001d0000000000000000000000000000001cffffffe3000000000000001d;
		6'b011110:	xpb = 256'h0000001e0000000000000000000000000000001dffffffe2000000000000001e;
		6'b011111:	xpb = 256'h0000001f0000000000000000000000000000001effffffe1000000000000001f;
		6'b100000:	xpb = 256'h000000200000000000000000000000000000001fffffffe00000000000000020;
		6'b100001:	xpb = 256'h0000002100000000000000000000000000000020ffffffdf0000000000000021;
		6'b100010:	xpb = 256'h0000002200000000000000000000000000000021ffffffde0000000000000022;
		6'b100011:	xpb = 256'h0000002300000000000000000000000000000022ffffffdd0000000000000023;
		6'b100100:	xpb = 256'h0000002400000000000000000000000000000023ffffffdc0000000000000024;
		6'b100101:	xpb = 256'h0000002500000000000000000000000000000024ffffffdb0000000000000025;
		6'b100110:	xpb = 256'h0000002600000000000000000000000000000025ffffffda0000000000000026;
		6'b100111:	xpb = 256'h0000002700000000000000000000000000000026ffffffd90000000000000027;
		6'b101000:	xpb = 256'h0000002800000000000000000000000000000027ffffffd80000000000000028;
		6'b101001:	xpb = 256'h0000002900000000000000000000000000000028ffffffd70000000000000029;
		6'b101010:	xpb = 256'h0000002a00000000000000000000000000000029ffffffd6000000000000002a;
		6'b101011:	xpb = 256'h0000002b0000000000000000000000000000002affffffd5000000000000002b;
		6'b101100:	xpb = 256'h0000002c0000000000000000000000000000002bffffffd4000000000000002c;
		6'b101101:	xpb = 256'h0000002d0000000000000000000000000000002cffffffd3000000000000002d;
		6'b101110:	xpb = 256'h0000002e0000000000000000000000000000002dffffffd2000000000000002e;
		6'b101111:	xpb = 256'h0000002f0000000000000000000000000000002effffffd1000000000000002f;
		6'b110000:	xpb = 256'h000000300000000000000000000000000000002fffffffd00000000000000030;
		6'b110001:	xpb = 256'h0000003100000000000000000000000000000030ffffffcf0000000000000031;
		6'b110010:	xpb = 256'h0000003200000000000000000000000000000031ffffffce0000000000000032;
		6'b110011:	xpb = 256'h0000003300000000000000000000000000000032ffffffcd0000000000000033;
		6'b110100:	xpb = 256'h0000003400000000000000000000000000000033ffffffcc0000000000000034;
		6'b110101:	xpb = 256'h0000003500000000000000000000000000000034ffffffcb0000000000000035;
		6'b110110:	xpb = 256'h0000003600000000000000000000000000000035ffffffca0000000000000036;
		6'b110111:	xpb = 256'h0000003700000000000000000000000000000036ffffffc90000000000000037;
		6'b111000:	xpb = 256'h0000003800000000000000000000000000000037ffffffc80000000000000038;
		6'b111001:	xpb = 256'h0000003900000000000000000000000000000038ffffffc70000000000000039;
		6'b111010:	xpb = 256'h0000003a00000000000000000000000000000039ffffffc6000000000000003a;
		6'b111011:	xpb = 256'h0000003b0000000000000000000000000000003affffffc5000000000000003b;
		6'b111100:	xpb = 256'h0000003c0000000000000000000000000000003bffffffc4000000000000003c;
		6'b111101:	xpb = 256'h0000003d0000000000000000000000000000003cffffffc3000000000000003d;
		6'b111110:	xpb = 256'h0000003e0000000000000000000000000000003dffffffc2000000000000003e;
		6'b111111:	xpb = 256'h0000003f0000000000000000000000000000003effffffc1000000000000003f;
	endcase
end
endmodule